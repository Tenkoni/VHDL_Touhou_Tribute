-- ****************************************************
--                    Proyecto Final   
-- ****************************************************
-- Integrantes:
--   Garrido Lopez Luis Enrique
--   Miramonte Sarabia Luis Enrique
--   Ortiz Figueroa Maria Fernanda
-- ****************************************************

-- ****************************************************
--        Modulo para dibujar el inicio del juego
-- ****************************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package start is
	procedure background_start(		
		-- xcur y ycur son los valores actuales del cursor, 
		-- es decir, las coordenadas del pixel que se está dibujando, 
		-- xpos y ypos son las coordenadas desde donde se empieza a dibujar
		signal xcur, ycur: in integer; 
		-- Los colores que tendrá el objeto dibujado, colores por pixel, 
		-- se pusieron en 12 bits, lo que nos da 4096 colores RRRRGGGGBBBB
		signal rgb: out std_logic_vector(11 downto 0); 
		-- Bandera que marca si se dibujara o no
		signal draw: out std_logic
	); 
end start;

package body start is 
	procedure background_start(
		-- Se declaran las variables auxiliares para manejar 
		-- los respectivos parametros del procedimiento
		signal xcur, ycur: in integer;
		signal rgb: out std_logic_vector(11 downto 0);
		signal draw: out std_logic) is
		
		-- Variable auxiliar para saber posición del dibujo el pixel
		variable pos_dx: integer := 0;
		variable pos_dy: integer := 0;
		
		-- Matriz para letrero
		type letrero is array (21 downto 0) of std_logic_vector(145 downto 0);
		constant touhou: letrero := (
			"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
			"10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010",
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"00001111111111111111111100000000001111111100000000001111000000000001111000011111000000000011111000000000011111111000000000011110000000000011110000",
			"00001111111111111111111100000000001111111100000000001111000000000001111000011111000000000011111000000000011111111000000000011110000000000011110000",
			"00001111111111111111111100000000110000000011000000001111000000000001111000011111000000000011111000000001100000000110000000011110000000000011110000",
			"00001111111111111111111100000000110000000011000000001111000000000001111000011111000000000011111000000001100000000110000000011110000000000011110000",
			"00001111111111111111111100000011000000000000110000001111000000000001111000011111000000000011111000000110000000000001100000011110000000000011110000",
			"00000000000111111000000000000011000000000000110000001111000000000001111000011111000000000011111000000110000000000001100000011110000000000011110000",
			"00000000000111111000000000001100000000000000001100001111000000000001111000011111111111111111111000011000000000000000011000011110000000000011110000",
			"00000000000111111000000000001100000000000000001100001111000000000001111000011111111111111111111000011000000000000000011000011110000000000011110000",
			"00000000000111111000000000000011000000000000110000001111000000000001111000011111111111111111111000000110000000000001100000011110000000000011110000",
			"00000000000111111000000000000011000000000000110000001111000000000001111000011111000000000011111000000110000000000001100000011110000000000011110000",
			"00000000000111111000000000000000110000000011000000001111000000000001111000011111000000000011111000000001100000000110000000011110000000000011110000",
			"00000000000111111000000000000000110000000011000000000111000000000001110000011111000000000011111000000001100000000110000000001110000000000011100000",
			"00000000000111111000000000000000001111111100000000000011111111111111100000011111000000000011111000000000011111111000000000000111111111111111000000",
			"00000000000111111000000000000000001111111100000000000001111111111111000000011111000000000011111000000000011111111000000000000011111111111110000000",
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010",
			"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
		
		type dibujo is array (24 downto 0) of std_logic_vector(24 downto 0);
		constant fantasma: dibujo := (
			"0000000111110000000000000",
			"0000011000001100000000000",
			"0000100000000010000000000",
			"0001000000000001000000000",
			"0010000000000000100000000",
			"0100000000000000010000000",
			"0100000000000000010000000",
			"1000000000000000001000000",
			"1000011000011000001000000",
			"1000010000001000001000000",
			"1000011000011000001000000",
			"1000000000000000001000000",
			"1000000111100000001000000",
			"1011100000001110001000000",
			"1000010000010000001000000",
			"1000010000010000001000000",
			"1011100000001110000100100",
			"1000000000000000000011010",
			"0100000000000000000000001",
			"0100000000000000000000001",
			"0010000000000000000000010",
			"0001000000000000000000010",
			"0000100000000000000001100",
			"0000011000000000000110000",
			"0000000111111111111000000");
		
	begin 
		-- La siguientes lineas se encargan de dibujar diferentes rectangulos
		-- de manera vertical para presentar un diseño de inicio del juego
		if(xcur>160 and xcur<=160+33 and ycur>240+45 and ycur<=480+45) then 
			rgb<= x"f00";
			draw <= '1';
		elsif(xcur>160+34 and xcur<=160+67 and ycur>280+45 and ycur<=480+45) then 
			rgb<= x"f40";
			draw <= '1';
		elsif(xcur>160+68 and xcur<=160+101 and ycur>200+45 and ycur<=480+45) then 
			rgb<= x"f80";
			draw <= '1';
		elsif(xcur>160+102 and xcur<=160+135 and ycur>190+45 and ycur<=480+45) then 
			rgb<= x"fb0";
			draw <= '1';
		elsif(xcur>160+136 and xcur<=160+169 and ycur>300+45 and ycur<=480+45) then 
			rgb<= x"ff0";
			draw <= '1';
		elsif(xcur>160+170 and xcur<=160+203 and ycur>260+45 and ycur<=480+45) then 
			rgb<= x"bf0";
			draw <= '1';
		elsif(xcur>160+204 and xcur<=160+237 and ycur>230+45 and ycur<=480+45) then 
			rgb<= x"8f0";
			draw <= '1';
		elsif(xcur>160+238 and xcur<=160+271 and ycur>280+45 and ycur<=480+45) then 
			rgb<= x"4f0";
			draw <= '1';
		elsif(xcur>160+272 and xcur<=160+305 and ycur>320+45 and ycur<=480+45) then 
			rgb<= x"0f0";
			draw <= '1';
		elsif(xcur>160+306 and xcur<=160+339 and ycur>340+45 and ycur<=480+45) then 
			rgb<= x"0F0";
			draw <= '1';
		elsif(xcur>160+340 and xcur<=160+373 and ycur>300+45 and ycur<=480+45) then 
			rgb<= x"0f4";
			draw <= '1';
		elsif(xcur>160+374 and xcur<=160+407 and ycur>270+45 and ycur<=480+45) then 
			rgb<= x"0f8";
			draw <= '1';
		elsif(xcur>160+408 and xcur<=160+441 and ycur>250+45 and ycur<=480+45) then 
			rgb<= x"0fb";
			draw <= '1';
		elsif(xcur>160+442 and xcur<=160+475 and ycur>260+45 and ycur<=480+45) then 
			rgb<= x"0ff";
			draw <= '1';
		elsif(xcur>160+476 and xcur<=160+509 and ycur>240+45 and ycur<=480+45) then 
			rgb<= x"0bf";
			draw <= '1';
		elsif(xcur>160+510 and xcur<=160+543 and ycur>210+45 and ycur<=480+45) then 
			rgb<= x"08f";
			draw <= '1';
		elsif(xcur>160+544 and xcur<=160+577 and ycur>230+45 and ycur<=480+45) then 
			rgb<= x"04f";
			draw <= '1';
		elsif(xcur>160+578 and xcur<=160+611 and ycur>200+45 and ycur<=480+45) then 
			rgb<= x"00f";
			draw <= '1';
		elsif(xcur>160+612 and xcur<=160+645 and ycur>240+45 and ycur<=480+45) then 
			rgb<= x"40f";
			draw <= '1';
		elsif(xcur>160+646 and xcur<=160+680 and ycur>210+45 and ycur<=480+45) then 
			rgb<= x"70d";
			draw <= '1';
		-- Se dibuja el titulo del juego
		elsif(xcur>160+229 and xcur<=160+375 and ycur>100+45 and ycur<=122+45) then
			pos_dx := (((160+375)-xcur));
			pos_dy := (((122+45)-ycur));
			
			if (touhou(pos_dy)(pos_dx) = '1') then
				rgb <= x"fff";
				draw <= '1';
			else
				draw <= '0';
			end if;
		-- Se dibuja dibujito del juego
		elsif(xcur>160+385 and xcur<=160+410 and ycur>100+45 and ycur<=125+45) then
			pos_dx := (((160+410)-xcur));
			pos_dy := (((125+45)-ycur));
			
			if (fantasma(pos_dy)(pos_dx) = '1') then
				rgb <= x"fff";
				draw <= '1';
			else
				draw <= '0';
			end if;
		else
			draw <= '0';
		end if;
	end background_start;
end start;