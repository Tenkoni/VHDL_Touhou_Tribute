-- ****************************************************
--                    Proyecto Final   
-- ****************************************************
-- Integrantes:
--   Garrido Lopez Luis Enrique
--   Miramonte Sarabia Luis Enrique
--   Ortiz Figueroa Maria Fernanda
-- ****************************************************

-- ****************************************************
--        Modulo para dibujar al los personajes
-- ****************************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package sprite is
	procedure figure(		
		-- xcur y ycur son los valores actuales del cursor, 
		-- es decir, las coordenadas del pixel que se está dibujando, 
		-- xpos y ypos son las coordenadas desde donde se empieza a dibujar
		signal xcur, ycur, xpos, ypos: in integer; 
		-- Los colores que tendrá el objeto dibujado, colores por pixel, 
		-- se pusieron en 12 bits, lo que nos da 4096 colores RRRRGGGGBBBB
		signal rgb: out std_logic_vector(11 downto 0); 
		-- Bandera que marca si se dibujara o no
		signal draw: out std_logic;
		-- contador para sprite
		signal count_sprite : in integer;
		-- Verifica si se dibujo el sprite de personaje
		signal charac: out std_logic_vector(1 downto 0);
		-- Verifica animación del sprite
		signal animationsignal: std_logic_vector(3 downto 0)
	); 
end sprite;

package body sprite is 
	procedure figure(
		-- Se declaran las variables auxiliares para manejar 
		-- los respectivos parametros del procedimiento
		signal xcur, ycur, xpos, ypos: in integer;
		signal rgb: out std_logic_vector(11 downto 0);
		signal draw: out std_logic;
		signal count_sprite: in integer;
		signal charac: out std_logic_vector(1 downto 0);
		signal animationsignal: std_logic_vector(3 downto 0)) is
		
		-- Variable auxiliar para saber posición del dibujo el pixel
		variable pos_dx: integer := 0;
		variable pos_dy: integer := 0;
		
		-- Matriz para manejar el sprite
		type rom_sprite is array (0 to 1174) of std_logic_vector(11 downto 0);
		-- Se define el mapa de bits para el sprite
		constant marisa1 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"384",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"242",x"223",x"334",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3A3",x"222",x"334",x"334",x"334",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"112",x"334",x"334",x"445",x"445",x"334",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3D3",x"000",x"112",x"233",x"334",x"445",x"556",x"556",x"374",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"242",x"112",x"112",x"222",x"334",x"334",x"445",x"556",x"223",x"373",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"343",x"434",x"334",x"223",x"011",x"222",x"223",x"334",x"345",x"223",x"222",x"343",x"3D3",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"000",x"534",x"857",x"656",x"334",x"111",x"111",x"112",x"223",x"445",x"334",x"545",x"545",x"112",x"242",x"3D3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"000",x"111",x"212",x"868",x"B8A",x"B9B",x"656",x"212",x"111",x"222",x"345",x"334",x"323",x"334",x"334",x"112",x"000",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"243",x"222",x"223",x"122",x"323",x"757",x"A8A",x"867",x"323",x"111",x"112",x"334",x"233",x"122",x"334",x"344",x"334",x"333",x"112",x"3A3",x"1F1",x"0F0",x"0F0",x"2F2",x"254",x"223",x"223",x"222",x"233",x"334",x"223",x"333",x"434",x"435",x"223",x"000",x"122",x"223",x"112",x"334",x"445",x"445",x"556",x"334",x"334",x"495",x"0F0",x"0F0",x"495",x"334",x"233",x"223",x"233",x"334",x"345",x"345",x"344",x"345",x"345",x"334",x"222",x"111",x"001",x"122",x"334",x"345",x"666",x"455",x"345",x"455",x"3E3",x"0F0",x"0F0",x"4D4",x"455",x"344",x"345",x"445",x"445",x"445",x"345",x"345",x"345",x"345",x"334",x"334",x"334",x"223",x"233",x"334",x"455",x"556",x"445",x"586",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4D4",x"5A6",x"455",x"445",x"445",x"445",x"445",x"445",x"334",x"334",x"233",x"223",x"223",x"223",x"334",x"445",x"586",x"4D5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"495",x"334",x"334",x"223",x"112",x"111",x"111",x"112",x"122",x"223",x"666",x"99A",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"222",x"777",x"777",x"655",x"666",x"776",x"877",x"988",x"CBB",x"FEE",x"FFF",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"5A5",x"222",x"111",x"888",x"FFF",x"FFF",x"FFE",x"FFF",x"FFF",x"DDC",x"CAA",x"FED",x"EFE",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"444",x"666",x"555",x"333",x"444",x"DCC",x"FED",x"A99",x"887",x"333",x"666",x"FFF",x"BFB",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"666",x"CCC",x"BBB",x"555",x"111",x"444",x"666",x"112",x"444",x"222",x"444",x"EEE",x"CFC",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"465",x"CCC",x"DDD",x"888",x"777",x"EEE",x"999",x"666",x"A99",x"FFF",x"CCC",x"555",x"AAA",x"EEE",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"373",x"666",x"CBB",x"AAA",x"777",x"DCC",x"EEE",x"DCD",x"FFF",x"EEE",x"DCC",x"FFF",x"999",x"666",x"BBB",x"BEB",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"322",x"777",x"AAA",x"777",x"898",x"FFF",x"CBB",x"AAA",x"AAA",x"999",x"DDD",x"FFF",x"999",x"444",x"666",x"999",x"7F7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"544",x"766",x"777",x"112",x"555",x"FEE",x"DCC",x"545",x"112",x"001",x"666",x"EEE",x"BBB",x"666",x"AAA",x"888",x"696",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"655",x"333",x"112",x"111",x"222",x"AAA",x"555",x"223",x"334",x"234",x"111",x"544",x"888",x"444",x"778",x"EDD",x"999",x"6C6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"223",x"223",x"122",x"223",x"233",x"223",x"222",x"223",x"344",x"334",x"334",x"233",x"112",x"001",x"112",x"222",x"677",x"777",x"999",x"4F4",x"0F0",x"0F0",x"0F0",x"1F1",x"364",x"222",x"223",x"334",x"344",x"345",x"334",x"334",x"344",x"345",x"334",x"334",x"223",x"223",x"112",x"111",x"112",x"112",x"111",x"223",x"575",x"3E3",x"0F0",x"0F0",x"666",x"222",x"223",x"334",x"445",x"445",x"345",x"345",x"445",x"445",x"345",x"334",x"334",x"223",x"000",x"000",x"000",x"112",x"223",x"223",x"112",x"111",x"242",x"2F2",x"0F0",x"111",x"233",x"334",x"444",x"445",x"445",x"445",x"445",x"345",x"345",x"344",x"344",x"334",x"334",x"111",x"000",x"000",x"111",x"333",x"334",x"223",x"112",x"111",x"242",x"2F2",x"666",x"233",x"334",x"344",x"445",x"445",x"344",x"334",x"334",x"344",x"445",x"445",x"344",x"334",x"223",x"001",x"000",x"112",x"334",x"445",x"334",x"112",x"445",x"555",x"555",x"CCC",x"556",x"334",x"334",x"445",x"334",x"222",x"222",x"223",x"334",x"445",x"556",x"445",x"334",x"334",x"112",x"000",x"112",x"334",x"334",x"233",x"445",x"BBC",x"CDC",x"2F2",x"EEE",x"BBC",x"667",x"233",x"122",x"111",x"111",x"111",x"223",x"334",x"556",x"566",x"556",x"344",x"334",x"223",x"001",x"222",x"334",x"334",x"445",x"BBC",x"CFC",x"4F4",x"0F0",x"3F3",x"BFB",x"BBB",x"777",x"111",x"000",x"000",x"000",x"111",x"223",x"445",x"556",x"445",x"334",x"234",x"223",x"111",x"223",x"223",x"555",x"BBB",x"CEC",x"3F3",x"0F0",x"0F0",x"0F0",x"2F2",x"EDD",x"EEE",x"778",x"000",x"000",x"000",x"000",x"667",x"AAA",x"AAA",x"9AA",x"999",x"778",x"556",x"222",x"112",x"566",x"CCC",x"AFA",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6F6",x"AFA",x"DCC",x"777",x"655",x"666",x"667",x"AAA",x"BBB",x"999",x"BCC",x"BBB",x"FFF",x"EEE",x"99A",x"889",x"DDE",x"9F9",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"7F7",x"8F8",x"CEC",x"FFF",x"777",x"111",x"211",x"421",x"111",x"221",x"BBB",x"BBB",x"BBB",x"CBB",x"8F8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F4",x"9A8",x"111",x"311",x"632",x"B64",x"632",x"211",x"211",x"110",x"363",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F3",x"352",x"632",x"843",x"D75",x"A64",x"742",x"321",x"100",x"3D3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"742",x"953",x"D75",x"D75",x"A54",x"532",x"110",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"842",x"953",x"C64",x"C65",x"B64",x"531",x"373",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3D3",x"632",x"953",x"A64",x"B64",x"953",x"421",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"674",x"953",x"A63",x"853",x"863",x"4E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"863",x"853",x"742",x"4E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E4",x"963",x"7B5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F3",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa2 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"373",x"343",x"586",x"5C5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3A4",x"223",x"445",x"445",x"556",x"474",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"111",x"345",x"445",x"445",x"666",x"445",x"474",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"122",x"223",x"445",x"445",x"445",x"445",x"344",x"223",x"373",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"122",x"334",x"333",x"334",x"344",x"345",x"334",x"334",x"111",x"373",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"3A4",x"112",x"334",x"234",x"223",x"223",x"334",x"334",x"334",x"334",x"222",x"323",x"233",x"3D3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"242",x"111",x"545",x"656",x"445",x"223",x"122",x"334",x"334",x"334",x"334",x"434",x"434",x"112",x"001",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"222",x"222",x"111",x"534",x"978",x"979",x"878",x"434",x"223",x"334",x"334",x"334",x"222",x"223",x"223",x"122",x"112",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"223",x"334",x"334",x"234",x"223",x"545",x"979",x"B9A",x"868",x"323",x"111",x"223",x"334",x"111",x"223",x"334",x"334",x"233",x"343",x"4C5",x"2F2",x"0F0",x"0F0",x"3E3",x"223",x"334",x"334",x"334",x"334",x"345",x"334",x"334",x"333",x"111",x"000",x"000",x"000",x"000",x"111",x"223",x"344",x"445",x"445",x"345",x"334",x"586",x"1F1",x"1F1",x"475",x"334",x"334",x"334",x"334",x"345",x"445",x"445",x"334",x"334",x"112",x"001",x"111",x"000",x"111",x"223",x"223",x"345",x"556",x"445",x"445",x"586",x"2F2",x"0F0",x"0F0",x"2F2",x"3E4",x"4C5",x"575",x"445",x"445",x"445",x"445",x"666",x"778",x"445",x"223",x"122",x"112",x"223",x"223",x"233",x"445",x"556",x"575",x"4D5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4D4",x"575",x"344",x"445",x"555",x"666",x"667",x"455",x"334",x"223",x"122",x"122",x"234",x"495",x"4D4",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C5",x"334",x"545",x"888",x"555",x"111",x"112",x"223",x"223",x"444",x"777",x"999",x"7C7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"474",x"334",x"777",x"FED",x"FED",x"AA9",x"887",x"A99",x"BBB",x"EDC",x"FFE",x"DFC",x"BFA",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"484",x"334",x"122",x"434",x"DCB",x"FFE",x"FFF",x"FFF",x"FFF",x"CCB",x"BBA",x"FFE",x"9F8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"223",x"777",x"888",x"444",x"544",x"DCB",x"DDD",x"DDD",x"AAA",x"332",x"666",x"BBB",x"8F8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"344",x"BBB",x"EEE",x"888",x"333",x"555",x"334",x"444",x"555",x"333",x"333",x"999",x"BEC",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"677",x"DDD",x"999",x"777",x"FFF",x"BBB",x"666",x"888",x"EEE",x"FFF",x"666",x"666",x"EEE",x"8F8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E4",x"888",x"AAA",x"555",x"CCC",x"EEE",x"BBB",x"FFF",x"FFF",x"A99",x"DCD",x"FEE",x"777",x"CCC",x"CDD",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"7B7",x"AAA",x"444",x"655",x"DDD",x"BAA",x"766",x"AAA",x"BAA",x"888",x"BAA",x"EEE",x"999",x"777",x"999",x"8D8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"888",x"556",x"111",x"444",x"BAB",x"CCC",x"777",x"000",x"111",x"777",x"BAA",x"CCC",x"555",x"555",x"889",x"676",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"555",x"444",x"223",x"223",x"222",x"666",x"888",x"223",x"000",x"000",x"000",x"222",x"444",x"444",x"334",x"CCC",x"BBB",x"8A9",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4A4",x"233",x"223",x"223",x"334",x"223",x"223",x"334",x"223",x"111",x"000",x"000",x"000",x"000",x"000",x"001",x"555",x"AAA",x"667",x"696",x"2F2",x"0F0",x"0F0",x"0F0",x"3E3",x"233",x"223",x"223",x"334",x"445",x"345",x"334",x"345",x"344",x"223",x"000",x"000",x"000",x"000",x"000",x"111",x"222",x"223",x"233",x"223",x"484",x"0F0",x"0F0",x"2F2",x"343",x"223",x"223",x"334",x"334",x"223",x"334",x"345",x"445",x"345",x"334",x"112",x"000",x"000",x"000",x"001",x"222",x"334",x"333",x"233",x"333",x"223",x"6C6",x"5F5",x"777",x"223",x"223",x"223",x"223",x"122",x"001",x"223",x"445",x"556",x"445",x"334",x"223",x"111",x"000",x"000",x"111",x"333",x"334",x"334",x"233",x"223",x"223",x"777",x"FFF",x"666",x"223",x"122",x"001",x"000",x"000",x"000",x"223",x"334",x"566",x"556",x"334",x"334",x"223",x"112",x"001",x"222",x"334",x"445",x"334",x"223",x"112",x"445",x"AAA",x"CCC",x"DDD",x"556",x"001",x"000",x"000",x"000",x"000",x"223",x"334",x"667",x"777",x"345",x"445",x"334",x"233",x"223",x"333",x"344",x"445",x"334",x"112",x"000",x"667",x"8B8",x"1F1",x"CCC",x"CCC",x"666",x"000",x"000",x"000",x"000",x"222",x"334",x"556",x"788",x"455",x"344",x"345",x"334",x"334",x"334",x"445",x"334",x"223",x"222",x"666",x"CDC",x"5F5",x"0F0",x"3F3",x"9E9",x"BBB",x"223",x"001",x"111",x"000",x"000",x"223",x"455",x"667",x"556",x"445",x"334",x"334",x"334",x"334",x"334",x"334",x"445",x"667",x"9CA",x"2F2",x"0F0",x"0F0",x"0F0",x"2F2",x"CCC",x"AAB",x"555",x"212",x"000",x"000",x"122",x"334",x"556",x"556",x"666",x"778",x"455",x"334",x"778",x"778",x"667",x"DDD",x"ADA",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6F6",x"9E9",x"ADA",x"AAA",x"777",x"667",x"999",x"889",x"9AA",x"889",x"788",x"899",x"455",x"222",x"999",x"BFB",x"8B9",x"BFC",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"9E9",x"9D9",x"EEE",x"DDD",x"777",x"999",x"999",x"A76",x"642",x"422",x"110",x"494",x"0F0",x"1F1",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6B6",x"222",x"311",x"421",x"632",x"C64",x"A53",x"632",x"321",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"252",x"632",x"843",x"A54",x"C65",x"C65",x"743",x"421",x"4A4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D3",x"632",x"953",x"B64",x"C65",x"D75",x"843",x"421",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"674",x"953",x"C64",x"C65",x"D65",x"843",x"452",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E3",x"843",x"A54",x"C64",x"D65",x"742",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"8A4",x"953",x"A53",x"B64",x"563",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"8A5",x"953",x"A53",x"5D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"8B5",x"A85",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"3F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa3 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"2F2",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"465",x"556",x"575",x"4E4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"222",x"334",x"445",x"666",x"455",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"233",x"334",x"345",x"334",x"556",x"445",x"343",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"223",x"334",x"333",x"334",x"455",x"556",x"334",x"484",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"111",x"234",x"223",x"111",x"334",x"344",x"445",x"334",x"233",x"4D5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"111",x"222",x"234",x"223",x"000",x"223",x"334",x"334",x"334",x"233",x"323",x"595",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"323",x"645",x"767",x"868",x"545",x"323",x"212",x"223",x"334",x"334",x"233",x"333",x"323",x"121",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4C5",x"234",x"334",x"656",x"868",x"DAC",x"C9B",x"968",x"534",x"212",x"223",x"334",x"334",x"222",x"212",x"222",x"222",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"354",x"223",x"234",x"233",x"334",x"556",x"767",x"768",x"445",x"323",x"211",x"001",x"112",x"223",x"223",x"122",x"334",x"334",x"233",x"4C5",x"0F0",x"0F0",x"0F0",x"4D4",x"111",x"223",x"234",x"334",x"334",x"334",x"334",x"334",x"334",x"233",x"112",x"000",x"000",x"000",x"000",x"112",x"223",x"334",x"445",x"445",x"344",x"3E3",x"0F0",x"0F0",x"3E4",x"354",x"233",x"334",x"334",x"334",x"334",x"233",x"334",x"344",x"445",x"334",x"122",x"111",x"111",x"112",x"223",x"334",x"556",x"455",x"455",x"4D4",x"1F1",x"0F0",x"0F0",x"0F0",x"2F2",x"5B5",x"344",x"334",x"223",x"111",x"001",x"122",x"334",x"445",x"445",x"334",x"223",x"223",x"223",x"234",x"344",x"475",x"4C5",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4A4",x"000",x"000",x"000",x"112",x"445",x"656",x"666",x"555",x"445",x"334",x"223",x"556",x"7C7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"112",x"333",x"777",x"AAA",x"DCB",x"DDC",x"EDD",x"DDC",x"DCB",x"BBB",x"EDD",x"EFD",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"345",x"888",x"EDD",x"FFF",x"FED",x"EDC",x"FFF",x"FFE",x"FFE",x"FEE",x"EED",x"CFC",x"8F7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"001",x"111",x"444",x"BBB",x"FFF",x"DDD",x"556",x"DDD",x"DDC",x"BAA",x"FED",x"AF9",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"232",x"333",x"766",x"566",x"222",x"998",x"CCC",x"112",x"444",x"333",x"443",x"DCC",x"9E9",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"444",x"888",x"FFF",x"999",x"000",x"000",x"434",x"333",x"777",x"777",x"555",x"888",x"DED",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"555",x"BBB",x"BBB",x"988",x"BBB",x"999",x"666",x"BBB",x"FFF",x"FFF",x"DDD",x"AAA",x"EFF",x"DFD",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"BBB",x"BAA",x"A99",x"EDD",x"EDD",x"CCB",x"FFF",x"FFF",x"CCC",x"CCC",x"FFF",x"CBB",x"CCC",x"FFF",x"7F7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"9B9",x"FFF",x"988",x"988",x"DDD",x"BBB",x"998",x"999",x"888",x"433",x"BAA",x"DDD",x"BAA",x"988",x"CCC",x"BFB",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"888",x"988",x"544",x"333",x"A99",x"CCC",x"CBB",x"222",x"000",x"000",x"444",x"999",x"877",x"988",x"AAA",x"DDD",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"575",x"434",x"111",x"000",x"000",x"333",x"888",x"989",x"334",x"223",x"111",x"000",x"001",x"001",x"223",x"BAB",x"EEE",x"EFE",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"223",x"111",x"000",x"000",x"000",x"000",x"334",x"667",x"445",x"334",x"234",x"223",x"223",x"223",x"112",x"112",x"778",x"999",x"8C8",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"343",x"111",x"000",x"000",x"000",x"111",x"233",x"334",x"334",x"445",x"345",x"344",x"334",x"334",x"334",x"334",x"223",x"112",x"112",x"223",x"595",x"2F2",x"1F1",x"494",x"223",x"122",x"000",x"000",x"000",x"111",x"233",x"334",x"334",x"445",x"445",x"445",x"445",x"445",x"345",x"445",x"445",x"445",x"334",x"223",x"223",x"233",x"444",x"BBB",x"112",x"223",x"111",x"000",x"000",x"112",x"233",x"334",x"334",x"445",x"455",x"445",x"445",x"445",x"445",x"344",x"334",x"344",x"445",x"334",x"334",x"223",x"223",x"344",x"DDD",x"444",x"112",x"000",x"112",x"222",x"334",x"334",x"334",x"345",x"445",x"556",x"445",x"445",x"445",x"445",x"334",x"233",x"112",x"112",x"233",x"334",x"223",x"334",x"AAA",x"FFF",x"A99",x"112",x"112",x"234",x"334",x"334",x"334",x"345",x"445",x"556",x"556",x"455",x"445",x"445",x"445",x"334",x"233",x"111",x"000",x"111",x"122",x"445",x"AAA",x"DDD",x"FEE",x"BBB",x"778",x"223",x"334",x"334",x"334",x"334",x"445",x"455",x"556",x"556",x"455",x"445",x"445",x"345",x"334",x"223",x"112",x"000",x"000",x"000",x"889",x"AFA",x"2F2",x"4F4",x"DFD",x"DCC",x"667",x"223",x"234",x"334",x"334",x"345",x"445",x"556",x"667",x"9AA",x"778",x"445",x"334",x"889",x"888",x"334",x"000",x"000",x"555",x"BBB",x"7E7",x"0F0",x"0F0",x"1F1",x"8E8",x"CCC",x"889",x"445",x"234",x"234",x"334",x"667",x"888",x"988",x"CA9",x"B99",x"889",x"899",x"9AA",x"AAA",x"BBB",x"888",x"888",x"9AA",x"AB9",x"5F5",x"0F0",x"0F0",x"0F0",x"1F1",x"DFD",x"FFF",x"BBB",x"889",x"888",x"999",x"DDD",x"A88",x"732",x"832",x"954",x"CAA",x"888",x"000",x"211",x"888",x"888",x"777",x"5C5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4F4",x"1F1",x"6F6",x"8F8",x"6F6",x"9C8",x"522",x"843",x"943",x"B54",x"743",x"100",x"100",x"110",x"000",x"121",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5D5",x"410",x"A53",x"B54",x"C64",x"843",x"421",x"211",x"210",x"242",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5B4",x"311",x"A53",x"C64",x"C64",x"A54",x"843",x"421",x"210",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"311",x"842",x"A54",x"C64",x"B54",x"843",x"421",x"4A3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"342",x"632",x"843",x"B54",x"B54",x"843",x"342",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"521",x"732",x"A53",x"B54",x"843",x"4A4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6D4",x"631",x"842",x"A54",x"753",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"6D4",x"974",x"A53",x"6D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F3",x"9A5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa4 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"373",x"343",x"343",x"495",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"373",x"334",x"345",x"334",x"445",x"343",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"343",x"334",x"445",x"345",x"556",x"445",x"223",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"334",x"334",x"334",x"334",x"445",x"556",x"334",x"243",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"222",x"334",x"223",x"233",x"334",x"334",x"445",x"344",x"223",x"494",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"001",x"233",x"344",x"334",x"223",x"223",x"334",x"334",x"334",x"334",x"333",x"474",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"232",x"323",x"545",x"445",x"334",x"234",x"223",x"112",x"223",x"334",x"334",x"334",x"323",x"112",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4D4",x"243",x"223",x"223",x"656",x"978",x"979",x"A89",x"756",x"433",x"112",x"223",x"334",x"233",x"111",x"223",x"223",x"4C5",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4D4",x"374",x"223",x"233",x"334",x"334",x"445",x"656",x"767",x"656",x"434",x"323",x"111",x"001",x"223",x"223",x"000",x"222",x"334",x"334",x"5A5",x"2F2",x"0F0",x"1F1",x"495",x"223",x"233",x"234",x"334",x"334",x"334",x"334",x"334",x"334",x"234",x"233",x"122",x"000",x"000",x"000",x"000",x"111",x"334",x"334",x"345",x"344",x"788",x"0F0",x"0F0",x"2F2",x"474",x"233",x"334",x"334",x"223",x"223",x"334",x"445",x"445",x"445",x"334",x"334",x"223",x"111",x"112",x"223",x"334",x"445",x"475",x"596",x"4D4",x"1F1",x"0F0",x"0F0",x"0F0",x"1F1",x"4A5",x"234",x"222",x"001",x"111",x"223",x"334",x"555",x"556",x"445",x"334",x"334",x"233",x"223",x"334",x"556",x"4E4",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4A5",x"001",x"000",x"000",x"111",x"223",x"334",x"444",x"445",x"334",x"334",x"334",x"445",x"667",x"989",x"7E7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"252",x"222",x"223",x"112",x"112",x"666",x"988",x"988",x"A99",x"A99",x"A99",x"BBA",x"EDD",x"DFC",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"223",x"122",x"111",x"766",x"FFE",x"FFE",x"DCB",x"DCC",x"FFE",x"FED",x"CFC",x"2F2",x"7F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"494",x"111",x"011",x"777",x"DCB",x"EDC",x"FFF",x"CCB",x"333",x"BBA",x"FFE",x"AF9",x"0F0",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E4",x"AAA",x"888",x"445",x"444",x"BAA",x"FED",x"BBA",x"666",x"000",x"444",x"AAA",x"7E7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6A6",x"FFF",x"DDD",x"777",x"444",x"444",x"666",x"112",x"556",x"556",x"333",x"665",x"CEC",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"777",x"DDD",x"877",x"655",x"EEE",x"CCC",x"556",x"777",x"CCC",x"DDD",x"BBB",x"777",x"AAA",x"9F9",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"484",x"989",x"888",x"433",x"999",x"CBB",x"BAA",x"FFF",x"CCC",x"777",x"AAA",x"EEE",x"999",x"766",x"CDC",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"565",x"AAA",x"544",x"333",x"AAA",x"BBB",x"888",x"999",x"666",x"333",x"A99",x"EDD",x"888",x"555",x"999",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"877",x"999",x"111",x"333",x"BAA",x"CBB",x"877",x"111",x"000",x"111",x"444",x"988",x"AAA",x"988",x"766",x"CFC",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"343",x"222",x"111",x"001",x"111",x"988",x"988",x"333",x"223",x"223",x"223",x"223",x"223",x"323",x"333",x"233",x"AAA",x"BFB",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"353",x"112",x"122",x"112",x"000",x"000",x"444",x"333",x"222",x"334",x"334",x"334",x"233",x"223",x"223",x"223",x"112",x"333",x"898",x"1F1",x"0F0",x"0F0",x"1F1",x"4A4",x"222",x"233",x"223",x"122",x"000",x"000",x"000",x"111",x"223",x"334",x"445",x"445",x"334",x"334",x"334",x"334",x"334",x"233",x"223",x"223",x"5A5",x"1F1",x"0F0",x"666",x"223",x"334",x"223",x"111",x"000",x"000",x"000",x"000",x"222",x"334",x"445",x"455",x"455",x"345",x"344",x"345",x"445",x"345",x"345",x"334",x"234",x"223",x"495",x"1F1",x"555",x"334",x"333",x"112",x"000",x"000",x"000",x"000",x"111",x"334",x"345",x"455",x"556",x"556",x"445",x"345",x"345",x"334",x"334",x"345",x"345",x"334",x"234",x"233",x"455",x"AAB",x"334",x"223",x"111",x"000",x"000",x"000",x"111",x"333",x"334",x"445",x"556",x"667",x"667",x"556",x"445",x"445",x"334",x"334",x"334",x"345",x"334",x"234",x"223",x"223",x"AAA",x"667",x"112",x"000",x"000",x"000",x"000",x"223",x"334",x"345",x"556",x"666",x"777",x"667",x"666",x"556",x"445",x"334",x"223",x"111",x"112",x"234",x"334",x"234",x"667",x"FFF",x"BBB",x"011",x"000",x"000",x"000",x"111",x"223",x"345",x"445",x"556",x"667",x"777",x"677",x"777",x"556",x"445",x"778",x"AAA",x"444",x"000",x"111",x"223",x"667",x"EEE",x"FFF",x"999",x"777",x"555",x"000",x"000",x"111",x"223",x"334",x"345",x"445",x"666",x"778",x"999",x"777",x"889",x"A9A",x"777",x"888",x"999",x"445",x"000",x"223",x"AAA",x"6F6",x"2F2",x"7D7",x"8F8",x"DCC",x"555",x"111",x"000",x"556",x"899",x"778",x"888",x"888",x"BBB",x"BBB",x"111",x"777",x"777",x"000",x"000",x"999",x"DDD",x"666",x"9B9",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"8F8",x"ADB",x"99A",x"666",x"A99",x"EEE",x"CCC",x"CCC",x"EEE",x"777",x"555",x"000",x"000",x"000",x"000",x"121",x"8C8",x"AFA",x"BEB",x"7F7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"7F7",x"EFE",x"5E5",x"1F1",x"2F2",x"544",x"655",x"210",x"310",x"000",x"110",x"210",x"110",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5F5",x"1F1",x"0F0",x"2F2",x"532",x"621",x"943",x"A54",x"522",x"421",x"320",x"362",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"732",x"943",x"C64",x"C65",x"B54",x"631",x"320",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"732",x"A53",x"C64",x"C64",x"B54",x"531",x"493",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"673",x"A53",x"B54",x"C54",x"C64",x"631",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"842",x"942",x"A53",x"B64",x"632",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"794",x"732",x"942",x"A53",x"743",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6D4",x"842",x"942",x"7A5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F3",x"974",x"8B5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F2",x"4F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa5 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"223",x"343",x"394",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"334",x"345",x"445",x"334",x"111",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"223",x"334",x"445",x"445",x"445",x"334",x"011",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"474",x"234",x"223",x"334",x"445",x"445",x"334",x"223",x"363",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"223",x"223",x"112",x"223",x"345",x"445",x"334",x"334",x"112",x"394",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"243",x"223",x"223",x"111",x"111",x"233",x"334",x"334",x"334",x"334",x"112",x"3A4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"343",x"434",x"334",x"334",x"223",x"111",x"112",x"223",x"334",x"334",x"334",x"223",x"112",x"495",x"4E4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"1F1",x"2F2",x"374",x"223",x"323",x"545",x"867",x"978",x"868",x"646",x"433",x"222",x"222",x"223",x"233",x"223",x"111",x"223",x"334",x"4C5",x"0F0",x"0F0",x"0F0",x"0F0",x"5B5",x"445",x"223",x"223",x"234",x"234",x"334",x"556",x"767",x"656",x"545",x"333",x"211",x"001",x"111",x"111",x"111",x"111",x"222",x"223",x"334",x"4C5",x"1F1",x"0F0",x"0F0",x"2F2",x"233",x"223",x"233",x"334",x"334",x"334",x"344",x"334",x"334",x"334",x"223",x"111",x"000",x"000",x"000",x"111",x"222",x"233",x"233",x"334",x"465",x"4E4",x"0F0",x"0F0",x"0F0",x"5A5",x"223",x"111",x"011",x"222",x"334",x"455",x"555",x"445",x"334",x"233",x"223",x"112",x"111",x"112",x"223",x"334",x"334",x"334",x"5B5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"494",x"111",x"000",x"000",x"222",x"344",x"445",x"445",x"334",x"334",x"223",x"112",x"122",x"223",x"234",x"234",x"344",x"4D5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4D4",x"253",x"000",x"111",x"122",x"334",x"334",x"334",x"334",x"233",x"445",x"887",x"988",x"999",x"DDD",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"3A4",x"222",x"222",x"334",x"444",x"555",x"888",x"BAA",x"FED",x"FDD",x"FED",x"FED",x"FFF",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"334",x"112",x"434",x"BA9",x"CBA",x"FED",x"FFE",x"FFE",x"FFE",x"FED",x"EEC",x"AF9",x"7F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"252",x"223",x"223",x"111",x"999",x"FFE",x"FED",x"FFF",x"CCB",x"AA9",x"FFD",x"9B8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4A4",x"444",x"445",x"444",x"000",x"222",x"BBA",x"888",x"988",x"555",x"332",x"CCB",x"ABA",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"333",x"DDD",x"DDD",x"545",x"333",x"222",x"111",x"333",x"444",x"333",x"111",x"AAA",x"DDD",x"6D6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"444",x"CCC",x"877",x"322",x"DDD",x"DDD",x"333",x"666",x"DDD",x"BBB",x"333",x"999",x"FFF",x"ACA",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"766",x"A9A",x"655",x"AAA",x"FFF",x"999",x"AAA",x"FFF",x"BBB",x"888",x"999",x"555",x"BBB",x"AAA",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"555",x"877",x"555",x"222",x"BBB",x"DDD",x"999",x"AAA",x"999",x"999",x"AAA",x"AAA",x"666",x"AAA",x"889",x"7E7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"888",x"444",x"111",x"000",x"444",x"BBB",x"CCC",x"BBB",x"111",x"111",x"888",x"988",x"444",x"999",x"AAA",x"999",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"766",x"555",x"112",x"222",x"222",x"111",x"001",x"444",x"889",x"445",x"000",x"111",x"333",x"222",x"111",x"111",x"555",x"999",x"2F2",x"0F0",x"0F0",x"2F2",x"5B5",x"484",x"464",x"223",x"112",x"223",x"334",x"223",x"222",x"111",x"000",x"222",x"223",x"000",x"111",x"334",x"345",x"223",x"112",x"001",x"111",x"474",x"2F2",x"0F0",x"CCD",x"334",x"112",x"223",x"223",x"223",x"334",x"334",x"223",x"334",x"223",x"000",x"000",x"000",x"001",x"223",x"334",x"445",x"445",x"334",x"222",x"112",x"223",x"343",x"3E3",x"AAA",x"223",x"223",x"223",x"223",x"334",x"445",x"334",x"334",x"233",x"111",x"000",x"000",x"000",x"222",x"334",x"445",x"455",x"555",x"445",x"334",x"223",x"223",x"233",x"444",x"AAA",x"122",x"223",x"223",x"334",x"445",x"445",x"334",x"334",x"112",x"000",x"000",x"000",x"112",x"223",x"334",x"556",x"667",x"667",x"445",x"334",x"223",x"112",x"223",x"334",x"778",x"223",x"223",x"334",x"334",x"334",x"334",x"223",x"112",x"111",x"000",x"000",x"112",x"223",x"334",x"445",x"556",x"667",x"667",x"889",x"767",x"666",x"223",x"000",x"222",x"CCD",x"556",x"223",x"334",x"334",x"223",x"222",x"111",x"000",x"000",x"001",x"112",x"223",x"334",x"345",x"445",x"667",x"878",x"DDD",x"DDD",x"BAA",x"FFF",x"AAA",x"666",x"666",x"CFC",x"ABA",x"677",x"223",x"233",x"222",x"001",x"000",x"000",x"112",x"223",x"334",x"334",x"334",x"334",x"445",x"DDD",x"BAA",x"888",x"222",x"333",x"AAA",x"A99",x"FFF",x"EEE",x"0F0",x"2F2",x"9F9",x"889",x"778",x"222",x"000",x"000",x"223",x"334",x"334",x"334",x"334",x"334",x"334",x"778",x"999",x"222",x"121",x"383",x"3E3",x"1F1",x"2F2",x"7F7",x"6F6",x"0F0",x"0F0",x"2F2",x"EEE",x"DDD",x"444",x"000",x"222",x"334",x"334",x"445",x"667",x"778",x"888",x"9AA",x"444",x"000",x"373",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"7F7",x"9D9",x"878",x"666",x"777",x"788",x"778",x"BBB",x"EEE",x"DDD",x"999",x"999",x"000",x"373",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"AFA",x"BEB",x"CBB",x"FFF",x"BAA",x"876",x"755",x"A76",x"732",x"100",x"000",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5F5",x"AFA",x"5E4",x"421",x"521",x"A43",x"B54",x"522",x"100",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"421",x"632",x"A54",x"C54",x"843",x"321",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"742",x"742",x"A53",x"C64",x"A54",x"532",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"773",x"953",x"943",x"B54",x"A54",x"532",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5A4",x"842",x"842",x"A53",x"943",x"663",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"421",x"632",x"842",x"732",x"5D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5A4",x"311",x"732",x"874",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"763",x"6C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F2",x"4F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa6 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"494",x"243",x"253",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"365",x"334",x"334",x"334",x"112",x"3A3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"334",x"445",x"445",x"445",x"344",x"111",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"233",x"333",x"334",x"445",x"445",x"445",x"223",x"122",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"234",x"223",x"233",x"334",x"445",x"445",x"334",x"223",x"223",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4A5",x"223",x"234",x"223",x"222",x"334",x"334",x"344",x"334",x"223",x"222",x"323",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"494",x"343",x"545",x"334",x"334",x"334",x"223",x"223",x"334",x"334",x"334",x"334",x"333",x"222",x"212",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"4D4",x"474",x"223",x"223",x"656",x"979",x"B8A",x"B8A",x"645",x"323",x"222",x"334",x"334",x"334",x"334",x"212",x"000",x"232",x"4D4",x"0F0",x"0F0",x"0F0",x"1F1",x"5B5",x"223",x"223",x"223",x"223",x"234",x"334",x"556",x"868",x"868",x"545",x"323",x"112",x"111",x"223",x"223",x"111",x"000",x"111",x"111",x"112",x"4D4",x"0F0",x"0F0",x"0F0",x"2F2",x"495",x"222",x"233",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"233",x"222",x"111",x"000",x"000",x"111",x"122",x"223",x"222",x"112",x"112",x"3E4",x"0F0",x"0F0",x"0F0",x"2F2",x"121",x"112",x"334",x"334",x"345",x"445",x"445",x"445",x"445",x"334",x"334",x"334",x"233",x"333",x"334",x"334",x"233",x"223",x"494",x"3E3",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"111",x"334",x"334",x"345",x"445",x"445",x"455",x"455",x"445",x"334",x"334",x"334",x"334",x"334",x"334",x"223",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"475",x"334",x"445",x"455",x"556",x"556",x"445",x"445",x"444",x"334",x"334",x"334",x"334",x"354",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"223",x"334",x"445",x"334",x"334",x"555",x"988",x"AAA",x"999",x"777",x"999",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3D3",x"222",x"223",x"223",x"877",x"998",x"DCB",x"FFD",x"FFE",x"FFF",x"FED",x"FDC",x"7F7",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"343",x"233",x"223",x"222",x"DCB",x"EDD",x"FFE",x"FFF",x"DDC",x"AAA",x"FFE",x"FDC",x"EDC",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"777",x"666",x"334",x"111",x"998",x"FFE",x"CBB",x"766",x"444",x"222",x"BAA",x"DCC",x"4F4",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"565",x"BBB",x"BBB",x"888",x"667",x"333",x"665",x"111",x"111",x"223",x"444",x"555",x"AAA",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"888",x"DDD",x"AAA",x"666",x"FFF",x"DDD",x"444",x"555",x"444",x"AAA",x"EEE",x"999",x"DDD",x"ACA",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"999",x"CCC",x"777",x"999",x"FFF",x"BBB",x"DDD",x"FFF",x"DDD",x"DDD",x"FFF",x"EEE",x"999",x"BBB",x"6C6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"222",x"777",x"888",x"333",x"DDD",x"EEE",x"999",x"988",x"888",x"A99",x"AAA",x"CCC",x"AAA",x"666",x"777",x"676",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5C5",x"444",x"888",x"334",x"001",x"666",x"CCC",x"AAA",x"222",x"000",x"222",x"888",x"777",x"222",x"777",x"AAA",x"999",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F3",x"565",x"888",x"666",x"111",x"112",x"111",x"444",x"777",x"111",x"112",x"222",x"444",x"555",x"112",x"222",x"778",x"CCC",x"3F3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"464",x"544",x"444",x"222",x"223",x"223",x"223",x"222",x"223",x"222",x"334",x"334",x"334",x"345",x"445",x"334",x"223",x"444",x"585",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"223",x"223",x"222",x"223",x"334",x"334",x"334",x"334",x"233",x"334",x"334",x"334",x"334",x"334",x"445",x"445",x"445",x"334",x"223",x"223",x"495",x"2F2",x"0F0",x"3E3",x"353",x"222",x"223",x"234",x"334",x"334",x"334",x"344",x"334",x"334",x"334",x"334",x"334",x"334",x"233",x"334",x"445",x"445",x"445",x"445",x"334",x"223",x"555",x"7A7",x"445",x"222",x"222",x"223",x"334",x"334",x"334",x"334",x"345",x"345",x"344",x"334",x"334",x"334",x"112",x"111",x"223",x"334",x"445",x"445",x"445",x"445",x"556",x"555",x"FFF",x"DDD",x"667",x"223",x"334",x"334",x"334",x"334",x"334",x"334",x"345",x"334",x"334",x"334",x"223",x"000",x"000",x"111",x"223",x"334",x"334",x"455",x"999",x"BBB",x"EEE",x"6F6",x"9E9",x"CCC",x"556",x"334",x"445",x"445",x"445",x"344",x"344",x"344",x"344",x"334",x"333",x"111",x"000",x"000",x"000",x"556",x"778",x"555",x"788",x"CFC",x"9D9",x"8F8",x"0F0",x"0F0",x"BFB",x"999",x"667",x"445",x"445",x"445",x"445",x"344",x"345",x"334",x"233",x"111",x"000",x"000",x"000",x"444",x"EEE",x"BCB",x"484",x"5E5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"5F5",x"DED",x"99A",x"667",x"556",x"445",x"345",x"345",x"334",x"112",x"000",x"000",x"001",x"556",x"888",x"CDC",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6F6",x"BDB",x"8E8",x"9B9",x"778",x"445",x"445",x"122",x"111",x"333",x"555",x"777",x"AAA",x"575",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F4",x"8A8",x"334",x"555",x"889",x"888",x"DDD",x"BBB",x"333",x"222",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"3E3",x"222",x"988",x"766",x"544",x"333",x"110",x"000",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"322",x"411",x"632",x"943",x"622",x"521",x"211",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"342",x"622",x"943",x"C64",x"A53",x"632",x"211",x"3A3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"473",x"622",x"A43",x"B54",x"B54",x"732",x"211",x"383",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"622",x"832",x"A54",x"B54",x"732",x"100",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"543",x"521",x"943",x"943",x"522",x"242",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6A4",x"411",x"622",x"732",x"521",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F2",x"442",x"421",x"522",x"583",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"553",x"663",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3F3",x"3F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa7 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"364",x"4A4",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"344",x"344",x"344",x"474",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"484",x"334",x"334",x"445",x"445",x"474",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"233",x"334",x"334",x"445",x"445",x"334",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"474",x"334",x"223",x"334",x"344",x"344",x"334",x"222",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"373",x"223",x"334",x"223",x"223",x"334",x"334",x"334",x"223",x"363",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"363",x"112",x"223",x"234",x"223",x"112",x"233",x"334",x"334",x"234",x"122",x"101",x"495",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"373",x"222",x"434",x"334",x"223",x"122",x"112",x"112",x"233",x"334",x"334",x"223",x"323",x"323",x"5B5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5B5",x"112",x"222",x"545",x"656",x"656",x"545",x"334",x"222",x"112",x"223",x"233",x"334",x"323",x"212",x"112",x"243",x"495",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"495",x"223",x"223",x"223",x"334",x"656",x"B8A",x"DAC",x"A8A",x"545",x"323",x"212",x"112",x"112",x"122",x"112",x"223",x"122",x"112",x"343",x"3E4",x"0F0",x"0F0",x"3E3",x"233",x"001",x"111",x"223",x"334",x"334",x"234",x"445",x"767",x"767",x"556",x"334",x"222",x"111",x"111",x"223",x"223",x"223",x"223",x"223",x"484",x"2F2",x"0F0",x"0F0",x"0F0",x"2F2",x"242",x"111",x"334",x"334",x"334",x"334",x"344",x"345",x"345",x"334",x"334",x"334",x"334",x"223",x"223",x"223",x"223",x"223",x"465",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"353",x"334",x"334",x"344",x"445",x"556",x"556",x"556",x"445",x"344",x"334",x"334",x"334",x"334",x"334",x"334",x"465",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"5B5",x"445",x"445",x"556",x"556",x"556",x"556",x"445",x"334",x"223",x"223",x"234",x"234",x"334",x"5A5",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"334",x"334",x"333",x"223",x"223",x"223",x"434",x"555",x"767",x"777",x"877",x"4D5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3D3",x"223",x"222",x"666",x"988",x"888",x"BA9",x"DCB",x"EDC",x"FEE",x"FFE",x"FED",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"444",x"334",x"112",x"BBA",x"FFF",x"FFF",x"FFF",x"FFF",x"EDD",x"998",x"FED",x"FED",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"464",x"BBB",x"999",x"555",x"544",x"FEE",x"FFE",x"BBA",x"AAA",x"445",x"211",x"CBB",x"CCB",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"666",x"EEE",x"FFF",x"AAA",x"000",x"777",x"777",x"111",x"222",x"000",x"000",x"555",x"BBA",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"444",x"CCC",x"DDD",x"666",x"555",x"999",x"222",x"223",x"222",x"555",x"222",x"444",x"DDD",x"DFD",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"242",x"555",x"999",x"666",x"777",x"EEE",x"CCC",x"BBB",x"FFF",x"BBB",x"CCC",x"BBB",x"333",x"999",x"DDD",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"383",x"444",x"CCC",x"333",x"222",x"CCC",x"BBB",x"666",x"777",x"AAA",x"888",x"AAA",x"EEE",x"444",x"444",x"777",x"6B6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"666",x"666",x"000",x"222",x"888",x"888",x"666",x"111",x"000",x"000",x"666",x"FFF",x"777",x"444",x"999",x"676",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"474",x"222",x"112",x"222",x"333",x"666",x"555",x"222",x"122",x"234",x"122",x"001",x"666",x"888",x"111",x"666",x"AAA",x"5A5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"494",x"112",x"223",x"334",x"334",x"334",x"333",x"223",x"223",x"334",x"334",x"334",x"233",x"112",x"222",x"223",x"112",x"222",x"223",x"494",x"4D4",x"2F2",x"0F0",x"4D4",x"233",x"112",x"334",x"334",x"334",x"334",x"234",x"233",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"233",x"223",x"223",x"233",x"223",x"353",x"2F2",x"344",x"111",x"334",x"334",x"334",x"233",x"223",x"223",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"445",x"445",x"445",x"344",x"334",x"233",x"333",x"333",x"223",x"444",x"233",x"122",x"334",x"334",x"223",x"223",x"222",x"223",x"334",x"445",x"445",x"344",x"334",x"223",x"334",x"345",x"445",x"445",x"445",x"445",x"334",x"233",x"333",x"777",x"889",x"666",x"223",x"334",x"223",x"111",x"000",x"222",x"334",x"445",x"455",x"445",x"445",x"334",x"112",x"223",x"334",x"445",x"445",x"445",x"334",x"234",x"334",x"788",x"BFB",x"7F7",x"DDD",x"888",x"233",x"111",x"000",x"001",x"223",x"344",x"445",x"556",x"555",x"445",x"334",x"111",x"111",x"223",x"334",x"334",x"334",x"445",x"778",x"999",x"ADA",x"2F2",x"0F0",x"FFF",x"888",x"333",x"000",x"000",x"223",x"344",x"445",x"445",x"555",x"555",x"445",x"334",x"111",x"000",x"111",x"112",x"122",x"445",x"999",x"EEE",x"CFC",x"0F0",x"0F0",x"0F0",x"2F2",x"8D8",x"666",x"111",x"555",x"CCD",x"999",x"777",x"99A",x"778",x"445",x"334",x"223",x"000",x"000",x"000",x"000",x"444",x"CCC",x"FFF",x"9E9",x"5F5",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"CFC",x"889",x"CCC",x"BFB",x"9D9",x"8E8",x"9F9",x"999",x"889",x"888",x"778",x"777",x"777",x"666",x"888",x"999",x"888",x"6E6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"7E7",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"BBB",x"FFF",x"AAA",x"666",x"BBB",x"666",x"888",x"343",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"483",x"322",x"788",x"555",x"100",x"000",x"100",x"000",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"473",x"621",x"310",x"521",x"632",x"210",x"311",x"242",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"473",x"943",x"843",x"C64",x"B54",x"522",x"411",x"373",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4A4",x"A53",x"B54",x"C65",x"C65",x"742",x"311",x"4B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"943",x"C64",x"C65",x"C65",x"842",x"332",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"843",x"A53",x"C64",x"C64",x"732",x"4A3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"5D4",x"832",x"A53",x"A54",x"643",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"874",x"942",x"843",x"5D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F3",x"843",x"874",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F3",x"6D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		constant marisa8 : rom_sprite := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"4C4",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"494",x"334",x"334",x"364",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B4",x"334",x"445",x"455",x"344",x"363",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"344",x"334",x"344",x"556",x"667",x"334",x"242",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4B5",x"334",x"233",x"334",x"445",x"556",x"445",x"233",x"363",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"233",x"334",x"223",x"223",x"334",x"345",x"445",x"334",x"222",x"383",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C4",x"343",x"223",x"234",x"233",x"223",x"223",x"334",x"334",x"334",x"233",x"111",x"495",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4C5",x"323",x"434",x"334",x"233",x"233",x"223",x"122",x"122",x"333",x"334",x"334",x"122",x"222",x"343",x"4C4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4A5",x"223",x"323",x"434",x"656",x"767",x"556",x"445",x"434",x"111",x"112",x"333",x"334",x"112",x"222",x"323",x"223",x"4A5",x"1F1",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"484",x"223",x"223",x"223",x"334",x"757",x"B9A",x"DAC",x"B8A",x"757",x"323",x"111",x"112",x"233",x"111",x"212",x"223",x"223",x"223",x"484",x"2F2",x"0F0",x"0F0",x"2F2",x"354",x"223",x"223",x"233",x"233",x"234",x"334",x"445",x"657",x"556",x"434",x"334",x"223",x"111",x"111",x"000",x"223",x"334",x"234",x"223",x"223",x"344",x"2F2",x"0F0",x"3E4",x"465",x"234",x"233",x"234",x"334",x"345",x"445",x"345",x"334",x"334",x"334",x"334",x"334",x"233",x"222",x"122",x"334",x"334",x"334",x"334",x"334",x"4D5",x"0F0",x"0F0",x"0F0",x"0F0",x"4D4",x"465",x"334",x"345",x"445",x"445",x"455",x"445",x"445",x"445",x"345",x"334",x"334",x"334",x"334",x"334",x"334",x"334",x"344",x"4D4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4C5",x"455",x"445",x"555",x"555",x"455",x"445",x"445",x"334",x"334",x"334",x"223",x"334",x"334",x"344",x"5A5",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"445",x"445",x"445",x"334",x"223",x"222",x"234",x"334",x"445",x"666",x"999",x"4E4",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"112",x"666",x"AAA",x"999",x"877",x"777",x"988",x"A99",x"CBB",x"EDC",x"DCB",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"454",x"111",x"110",x"888",x"BAA",x"DCC",x"EDD",x"FFF",x"FEE",x"CBA",x"988",x"777",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"AAA",x"999",x"555",x"211",x"333",x"DDD",x"BAA",x"AAA",x"666",x"000",x"888",x"BBB",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"464",x"CCC",x"FFF",x"AAA",x"555",x"555",x"445",x"001",x"111",x"000",x"111",x"BBB",x"FFF",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"222",x"BBB",x"AAA",x"333",x"CCC",x"DDD",x"999",x"666",x"CCC",x"CCC",x"888",x"999",x"DDD",x"DED",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4A4",x"666",x"888",x"333",x"777",x"DDD",x"999",x"FFF",x"FFF",x"888",x"999",x"CCC",x"444",x"AAA",x"CCC",x"6E6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"343",x"EEE",x"667",x"111",x"AAA",x"CCC",x"777",x"666",x"888",x"666",x"777",x"CCC",x"555",x"666",x"999",x"8B8",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"494",x"999",x"889",x"222",x"111",x"888",x"999",x"333",x"000",x"000",x"111",x"777",x"BBB",x"777",x"999",x"AAA",x"888",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"556",x"667",x"112",x"222",x"112",x"777",x"666",x"223",x"223",x"223",x"112",x"222",x"555",x"666",x"334",x"CCC",x"999",x"494",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4A4",x"334",x"222",x"223",x"334",x"222",x"223",x"233",x"334",x"445",x"445",x"334",x"223",x"222",x"223",x"122",x"223",x"455",x"454",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"343",x"223",x"223",x"334",x"334",x"334",x"334",x"345",x"445",x"345",x"445",x"344",x"334",x"334",x"334",x"223",x"222",x"112",x"222",x"222",x"384",x"2F2",x"0F0",x"2F2",x"223",x"223",x"223",x"233",x"334",x"445",x"445",x"445",x"345",x"334",x"334",x"445",x"345",x"334",x"334",x"334",x"334",x"334",x"223",x"223",x"222",x"222",x"343",x"3D4",x"999",x"223",x"223",x"223",x"334",x"345",x"445",x"334",x"334",x"334",x"233",x"334",x"445",x"445",x"445",x"334",x"334",x"334",x"334",x"334",x"233",x"223",x"222",x"222",x"334",x"999",x"334",x"223",x"233",x"334",x"445",x"344",x"334",x"223",x"222",x"122",x"334",x"344",x"445",x"445",x"445",x"345",x"334",x"334",x"334",x"334",x"223",x"333",x"777",x"AAA",x"EEE",x"788",x"223",x"233",x"334",x"345",x"334",x"223",x"112",x"000",x"111",x"334",x"445",x"445",x"455",x"555",x"455",x"445",x"334",x"334",x"233",x"334",x"778",x"DDD",x"FFF",x"8F8",x"DDD",x"778",x"233",x"334",x"334",x"223",x"112",x"000",x"001",x"112",x"334",x"445",x"445",x"555",x"556",x"556",x"445",x"445",x"334",x"445",x"999",x"DDD",x"8E8",x"1F1",x"0F0",x"9F9",x"CCC",x"99A",x"445",x"233",x"112",x"000",x"333",x"AAB",x"99A",x"667",x"345",x"445",x"555",x"556",x"556",x"445",x"334",x"666",x"AAA",x"BFB",x"7F7",x"0F0",x"0F0",x"0F0",x"1F1",x"DFD",x"FFF",x"AAA",x"334",x"333",x"666",x"889",x"BBB",x"898",x"666",x"999",x"777",x"455",x"445",x"455",x"556",x"778",x"BBB",x"CFC",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4F4",x"5F5",x"CDC",x"BBB",x"BBC",x"CCC",x"333",x"000",x"000",x"011",x"888",x"898",x"99A",x"999",x"778",x"BBC",x"CDC",x"7F7",x"6F6",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"6F6",x"ADA",x"DDD",x"AAA",x"000",x"111",x"210",x"411",x"210",x"111",x"899",x"999",x"8C8",x"7F7",x"4F4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"4F4",x"5F5",x"4B4",x"210",x"522",x"B54",x"842",x"411",x"100",x"111",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"422",x"732",x"C64",x"B54",x"A53",x"521",x"111",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1F1",x"442",x"832",x"B54",x"C64",x"C54",x"632",x"221",x"2F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"463",x"832",x"A43",x"C64",x"B54",x"622",x"352",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"483",x"732",x"942",x"A53",x"943",x"522",x"3E3",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2F2",x"643",x"732",x"832",x"732",x"6B4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E3",x"642",x"732",x"843",x"3F2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"3E3",x"643",x"894",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"4E4",x"4E4",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");

	begin 
		
		-- Se dibuja al personaje del juego con una ilución de movimiento
		if(xcur>xpos and xcur<=xpos+25 and ycur>ypos and ycur<=ypos+47) then 
			draw <= '1';
			if(count_sprite < 1175) then
				if(animationsignal = x"0") then
					if (marisa1(count_sprite) /= x"0F0") then
						rgb<= marisa1(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;
					
				if(animationsignal = x"1") then
					if (marisa2(count_sprite) /= x"0F0") then
						rgb<= marisa2(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;
					
				if(animationsignal = x"2") then
					if (marisa3(count_sprite) /= x"0F0") then
						rgb<= marisa3(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;

				if(animationsignal = x"3") then
					
					if (marisa4(count_sprite) /= x"0F0") then
						rgb<= marisa4(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;

				if(animationsignal = x"4") then
					if (marisa5(count_sprite) /= x"0F0") then
						rgb<= marisa5(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;
					
				if(animationsignal = x"5") then
					if (marisa6(count_sprite) /= x"0F0") then
						rgb<= marisa6(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;
					
				if(animationsignal = x"6") then
					if (marisa7(count_sprite) /= x"0F0") then
						rgb<= marisa7(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;

				if(animationsignal = x"7") then
					if (marisa8(count_sprite) /= x"0F0") then
						rgb<= marisa8(count_sprite);
						-- Tiene la función como un draw exclusivo para el personaje
						-- [01 dibujo] [00 no dibujo] [10 transparencia] [11 reset]
						charac <="01"; 
					else 
						charac <= "10";
					end if;
				end if;
					
				if(count_sprite = 1174) then
					charac <= "11";
				end if;
			end if;
   	else
			draw <= '0';
			charac <= "00";
		end if;
	end figure;
end sprite;