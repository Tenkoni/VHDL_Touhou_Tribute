-- ****************************************************
--                    Proyecto Final   
-- ****************************************************
-- Integrantes:
--   Garrido Lopez Luis Enrique
--   Miramonte Sarabia Luis Enrique
--   Ortiz Figueroa Maria Fernanda
-- ****************************************************

-- ****************************************************
--        Módulo para dibujar los fondos y datos
--         de cada uno de los diferentes niveles
-- ****************************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package background is
	procedure background_play(		
		-- xcur y ycur son los valores actuales del cursor, 
		-- es decir, las coordenadas del pixel que se está dibujando, 
		-- xpos y ypos son las coordenadas desde donde se empieza a dibujar
		signal xcur, ycur: in integer; 
		-- Los colores que tendrá el objeto dibujado, colores por pixel, 
		-- se pusieron en 12 bits, lo que nos da 4096 colores RRRRGGGGBBBB
		signal rgb: out std_logic_vector(11 downto 0);
		-- Nivel
		signal nivel: in integer;
		-- Vida
		signal life: in integer;
		-- Score
		signal sc_u,sc_d,sc_c,sc_m,sc_mm: in integer
	); 
end background;

package body background is 
	procedure background_play(
		-- Se declaran las variables auxiliares para manejar 
		-- los respectivos parametros del procedimiento
		signal xcur, ycur: in integer;
		signal rgb: out std_logic_vector(11 downto 0);
		signal nivel: in integer;
		signal life: in integer;
		signal sc_u,sc_d,sc_c,sc_m,sc_mm: in integer) is
		
		-- Variable auxiliar para saber posición del dibujo el pixel
		variable pos_dx: integer := 0;
		variable pos_dy: integer := 0;
		
		-- Variables auxiliares para pintar el fondo
		variable y: integer;
		variable x: integer;
		
		-- Variables auxiliares para verificar que es lo que se pinta
		variable ay: integer;
		variable ax: integer;
		variable ac: integer;
		variable ae: integer;
		variable al: integer;
		
		-- Matriz para manejar el controno de la zona de datos(nombre, vidas score)
		type rom_datos is array (9 downto 0) of std_logic_vector (9 downto 0);
		-- Se define el mapa de bits para el margen de los datos
		constant margen_h : rom_datos := ("1111111111",
												    "1111111111",
												    "0000110000",
												    "0001111000",
												    "0011001100",
												    "0110000110",
												    "1100000011",
												    "1000000001",
												    "1111111111",
												    "1111111111");
												  
		-- Se define el mapa de bits para el margen de los datos
		constant margen_v : rom_datos := ("1111000011",
												    "1101100011",
												    "1100110011",
												    "1100011011",
												    "1100001111",
												    "1100001111",
												    "1100011011",
												    "1100110011",
												    "1101100011",
												    "1111000011");
													 
		-- Matris para manejar numeros
		type rom_numero is array (0 to 14) of std_logic_vector(0 to 14);
		constant uno : rom_numero := ( "000000111000000",	
												 "000011111000000",
												 "000011111000000",
												 "001100111000000",
												 "001100111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "000000111000000",
												 "011111111111110",
												 "011111111111110");
		constant dos : rom_numero := ( "000011111111100",
												 "000110000000110",
												 "001100000000110",
												 "000000000000110",
												 "000000000000110",
												 "000000000000110",
												 "000000000001100",
												 "000000000110000",
												 "000000011000000",
												 "000001100000000",
												 "000110000000000",
												 "011000000000000",
												 "011000000000000",
												 "011111111111110",
												 "011111111111110");
		constant tres : rom_numero := ( "000111111111000",
												  "011111111111100",
												  "011000000000110",
												  "000000000000110",
												  "000000000000110",
												  "000000000000110",
												  "000000000111100",
												  "000000000111100",
												  "000000000000110",
												  "000000000000110",
												  "000000000000110",
												  "011000000000110",
												  "011111111111110",
												  "000111111111000",
												  "000011111110000");
		constant cuatro : rom_numero := ( "011000000000110",
													 "011000000000110",
													 "011000000000110",
													 "011000000000110",
													 "011000000000110",
													 "011000000000110",
													 "001111111111110",
													 "000111111111110",
													 "000000000000110",
													 "000000000000110",
													 "000000000000110",
													 "000000000000110",
													 "000000000000110",
													 "000000000000110",
													 "000000000000110");
		constant cinco : rom_numero := ( "011111111111110",
													"011111111111110",
													"011000000000000",
													"011000000000000",
													"011000000000000",
													"011000000000000",
													"011111111111000",
													"000111111111000",
													"000000000000110",
													"000000000000110",
													"011000000000110",
													"011000000000110",
													"000111111111100",
													"000111111111100",
													"000011111111000");
		constant seis : rom_numero := ( "000001111111000",
												  "001111111111100",
												  "001110000001100",
												  "011000000000000",
												  "011000000000000",
												  "011000000000000",
												  "011000000000000",
												  "011111111111110",
												  "011111111111110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "000111111111100",
												  "000111111111000",
												  "000011111110000");
		constant siete : rom_numero := ( "000111111111110",
													"000111111111110",
													"011000000000110",
													"011000000000110",
													"000000000000110",
													"000000000011100",
													"000000000011100",
													"000000001100000",
													"000000001100000",
													"000000001100000",
													"000000001100000",
													"000000001100000",
													"000000001100000",
													"000000001100000",
													"000000001100000");
		constant ocho : rom_numero := ( "000111111111000",
												  "000111111111000",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "000111111111000",
												  "000111111111000",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011111111111110",
												  "000111111111000");
		constant nueve : rom_numero := ( "000001111111110",
													"000011111111110",
													"000110000000110",
													"001100000000110",
													"001100000000110",
													"001100000000110",
													"000110000000110",
													"000011111111110",
													"000011111111110",
													"000000000000110",
													"000000000000110",
													"000000000000110",
													"000000000000110",
													"000000000000110",
													"000000000000110");
		constant cero : rom_numero := ( "000111111111000",
												  "001111111111100",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "011000000000110",
												  "001111111111100",
												  "000111111111000");
		
		-- Matriz para manejar letreros 
		type rom_letrero is array(0 to 14) of std_logic_vector(0 to 74);
		constant l_score : rom_letrero := ( "001111111111100000001111111110000111111111000000111111111000011111111111110",
														"001111111111100000011111111110011111111111110000111111111100011111111111110",
														"011000000000110000110000000000011000000000110011000000000110011000000000000",
														"011000000000110001110000000000011000000000110011000000000110011000000000000",
														"011000000000000011000000000000011000000000110011000000000110011000000000000",
														"011000000000000011000000000000011000000000110011000000000110011000000000000",
														"000111111111000011000000000000011000000000110011000000001100011111111110000",
														"000111111111000011000000000000011000000000110011111111110000011111111110000",
														"000000000000110011000000000000011000000000110011001100000000011000000000000",
														"000000000000110011000000000000011000000000110011001100000000011000000000000",
														"000000000000110011000000000000011000000000110011000011000000011000000000000",
														"001100000000110001110000000000011000000000110011000000111000011000000000000",
														"001100000000110000110000000000011000000000110011000000000110011000000000000",
														"001111111111100000011111111110011111111111110011000000000110011111111111110",
														"000011111110000000001111111110000111111111000011000000000110011111111111110");
		constant l_nivel : rom_letrero := ( "011110000000110011111111111110011000000000110011111111111110011000000000000",
														"011110000000110011111111111110011000000000110011111111111110011000000000000",
														"011111000000110000000111000000011000000000110011000000000000011000000000000",
														"011011000000110000000111000000011000000000110011000000000000011000000000000",
														"011001100000110000000111000000001100000001100011000000000000011000000000000",
														"011001100000110000000111000000001100000001100011000000000000011000000000000",
														"011000110000110000000111000000001100000001100011111111110000011000000000000",
														"011000110000110000000111000000001100000001100011111111110000011000000000000",
														"011000011000110000000111000000000111000111000011000000000000011000000000000",
														"011000011000110000000111000000000011000110000011000000000000011000000000000",
														"011000001100110000000111000000000011000110000011000000000000011000000000000",
														"011000001100110000000111000000000011000110000011000000000000011000000000000",
														"011000000110110000000111000000000001101100000011000000000000011000000000000",
														"011000000111110011111111111110000000111000000011111111111110011111111111110",
														"011000000011110011111111111110000000010000000011111111111110011111111111110");
		
		-- Matriz para manejar un diseño del fondo
		type rom_fondo is array (0 to 1919) of std_logic_vector(11 downto 0);
		-- Se define el mapa de bits para el piso del fondo
		constant piso1 : rom_fondo := ( x"834",x"834",x"733",x"843",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"834",x"834",x"733",x"733",x"833",x"744",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"200",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"000",x"000",x"000",x"000",x"834",x"833",x"843",x"743",x"743",x"744",x"000",x"100",x"C84",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C84",x"100",x"100",x"C84",x"E82",x"D82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D84",x"100",x"100",x"D83",x"E82",x"E82",x"E82",x"E82",x"E92",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C83",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"733",x"744",x"743",x"644",x"644",x"000",x"100",x"E82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F70",x"F80",x"F70",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F70",x"F70",x"F70",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"D82",x"100",x"000",x"000",x"000",x"000",x"000",x"733",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"200",x"200",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E83",x"100",x"100",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"000",x"000",x"000",x"744",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E81",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"E82",x"200",x"200",x"E82",x"F70",x"F80",x"F70",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"100",x"D82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"D82",x"200",x"000",x"000",x"000",x"000",x"000",x"843",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"E82",x"200",x"100",x"D84",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D84",x"100",x"100",x"D94",x"D82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D94",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"743",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"000",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"645",x"744",x"744",x"643",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"744",x"734",x"733",x"844",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"C83",x"E82",x"E82",x"E82",x"E82",x"E83",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D82",x"E82",x"E83",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C83",x"100",x"100",x"744",x"834",x"844",x"733",x"833",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E81",x"100",x"100",x"734",x"834",x"833",x"844",x"833",x"733",x"743",x"743",x"743",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"734",x"834",x"833",x"733",x"844",x"733",x"843",x"833",x"833",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"744",x"733",x"844",x"733",x"734",x"734",x"833",x"833",x"833",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"200",x"E82",x"F70",x"F80",x"F70",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"D81",x"100",x"000",x"744",x"844",x"733",x"743",x"734",x"734",x"734",x"834",x"834",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"E82",x"100",x"100",x"E82",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"000",x"644",x"734",x"744",x"743");
		constant piso2 : rom_fondo := ( x"834",x"834",x"733",x"843",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"834",x"834",x"733",x"733",x"833",x"744",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"200",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"200",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"000",x"000",x"000",x"000",x"834",x"833",x"843",x"743",x"743",x"744",x"000",x"100",x"C84",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C84",x"100",x"100",x"C84",x"E82",x"D82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D84",x"100",x"100",x"D83",x"E82",x"E82",x"E82",x"E82",x"E92",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E83",x"E83",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C83",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"733",x"744",x"743",x"644",x"644",x"000",x"100",x"E82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F70",x"F80",x"F70",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F81",x"F81",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F70",x"F70",x"F70",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"D82",x"100",x"000",x"000",x"000",x"000",x"000",x"733",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"200",x"200",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E83",x"100",x"100",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"000",x"000",x"000",x"744",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E81",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"E82",x"200",x"200",x"E82",x"F70",x"F80",x"F70",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"100",x"D82",x"F80",x"F80",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"D82",x"200",x"000",x"000",x"000",x"000",x"000",x"843",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"E82",x"200",x"100",x"D84",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D84",x"100",x"100",x"D94",x"D82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E81",x"E82",x"E82",x"D82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D94",x"100",x"000",x"000",x"000",x"000",x"000",x"833",x"743",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"000",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"645",x"744",x"744",x"643",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"200",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"100",x"000",x"000",x"744",x"734",x"733",x"844",x"833",x"744",x"000",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"C83",x"E82",x"E82",x"E82",x"E82",x"E83",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D82",x"E82",x"E83",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"D84",x"100",x"100",x"D84",x"E82",x"E82",x"E83",x"E82",x"E82",x"E82",x"E82",x"E81",x"E81",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"E82",x"C83",x"100",x"100",x"744",x"834",x"844",x"733",x"833",x"744",x"100",x"000",x"000",x"000",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"200",x"200",x"E82",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E81",x"100",x"100",x"734",x"834",x"833",x"844",x"833",x"733",x"743",x"743",x"743",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F70",x"F80",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"000",x"734",x"834",x"833",x"733",x"844",x"733",x"843",x"833",x"833",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F70",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F70",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"744",x"733",x"844",x"733",x"734",x"734",x"833",x"833",x"833",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"200",x"E82",x"F70",x"F80",x"F70",x"F80",x"F80",x"F80",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E81",x"F80",x"F70",x"F80",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"D81",x"100",x"000",x"744",x"844",x"733",x"743",x"734",x"734",x"734",x"834",x"834",x"744",x"000",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F70",x"F70",x"E82",x"100",x"100",x"E82",x"F70",x"F70",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"E82",x"100",x"100",x"E82",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F80",x"F70",x"E82",x"100",x"000",x"644",x"734",x"744",x"743");
		constant piso3 : rom_fondo := ( x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222");
		constant piso4 : rom_fondo := ( x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"FFF",x"FFF",x"333",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"333",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222",x"222");		
		
		-- Matriz para manejar un diseño del fondo
		type rom_cosas is array (0 to 623) of std_logic_vector(11 downto 0);
		-- Se define el mapa de bits para las flores del fondo
		constant flores : rom_cosas := ( x"00F",x"00F",x"00F",x"00C",x"FFF",x"FFF",x"00C",x"30B",x"C04",x"F00",x"C00",x"904",x"20B",x"00C",x"FFF",x"FFF",x"00C",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00E",x"00D",x"008",x"FFF",x"FFF",x"008",x"308",x"C14",x"E00",x"D00",x"A03",x"208",x"018",x"FFF",x"FFF",x"018",x"00C",x"00C",x"00D",x"00E",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00D",x"FFF",x"FFF",x"FF7",x"FF7",x"FFF",x"FEF",x"A01",x"D00",x"E00",x"C12",x"FEF",x"FFF",x"FF6",x"FF7",x"FFF",x"FFF",x"FFF",x"EEF",x"00D",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00B",x"EFF",x"FFB",x"EF5",x"FF6",x"FFC",x"FFE",x"820",x"910",x"B13",x"A24",x"FFE",x"FFB",x"FF6",x"FE5",x"FFC",x"FFE",x"FFD",x"FFF",x"109",x"10B",x"30B",x"30B",x"20B",x"20B",x"00F",x"01B",x"7BA",x"8C6",x"FFC",x"FFD",x"140",x"140",x"9B5",x"AA8",x"207",x"207",x"8B8",x"8C5",x"FFB",x"FFD",x"FFF",x"FFD",x"FE6",x"FF7",x"FFF",x"FEF",x"A15",x"C04",x"A04",x"904",x"00F",x"01A",x"6B9",x"7D5",x"DFD",x"EFE",x"140",x"050",x"7D5",x"7C9",x"01A",x"00A",x"9B9",x"AB5",x"FFD",x"FEF",x"FEF",x"FFF",x"FE7",x"EE7",x"FFF",x"FEF",x"C11",x"F00",x"D00",x"C00",x"00F",x"01A",x"7C9",x"6D4",x"7D5",x"7C6",x"140",x"040",x"6C4",x"7C8",x"01A",x"20B",x"713",x"910",x"C10",x"A14",x"308",x"109",x"FFF",x"FFF",x"018",x"208",x"A03",x"C00",x"E00",x"F00",x"20B",x"207",x"AA8",x"9B5",x"7C7",x"7C8",x"040",x"140",x"7C5",x"7B8",x"117",x"407",x"A03",x"D00",x"E00",x"C14",x"30B",x"00C",x"FFF",x"EFF",x"01C",x"10B",x"714",x"A11",x"C13",x"C04",x"C04",x"C13",x"C11",x"923",x"107",x"017",x"143",x"140",x"050",x"130",x"723",x"A03",x"D01",x"F00",x"F00",x"C04",x"30B",x"00B",x"134",x"134",x"00B",x"00B",x"334",x"322",x"307",x"30B",x"F00",x"F00",x"F00",x"C14",x"208",x"028",x"032",x"140",x"040",x"340",x"620",x"A10",x"D10",x"E01",x"C03",x"917",x"208",x"017",x"042",x"042",x"018",x"028",x"032",x"143",x"018",x"00B",x"C00",x"D00",x"F00",x"C12",x"423",x"033",x"141",x"140",x"140",x"140",x"9B5",x"CA5",x"A10",x"A03",x"508",x"108",x"8BB",x"7C8",x"050",x"141",x"032",x"143",x"041",x"041",x"143",x"134",x"904",x"A02",x"C12",x"A21",x"330",x"140",x"150",x"050",x"040",x"050",x"7D5",x"9C5",x"620",x"713",x"107",x"026",x"7C7",x"7D4",x"040",x"140",x"140",x"140",x"140",x"140",x"040",x"040",x"20B",x"208",x"423",x"330",x"240",x"050",x"7C5",x"6C5",x"6D5",x"7D5",x"6C4",x"7C5",x"240",x"230",x"8C8",x"7C8",x"6D5",x"6D4",x"AE6",x"AD5",x"AD5",x"BD6",x"AD5",x"AD7",x"140",x"040",x"00F",x"00C",x"137",x"143",x"040",x"050",x"7C4",x"7D4",x"7D4",x"6D4",x"7D4",x"7C5",x"040",x"050",x"7C4",x"6D4",x"6D4",x"7D4",x"AD4",x"BD4",x"BD5",x"BD5",x"BD5",x"AD7",x"140",x"040",x"00F",x"00E",x"00C",x"018",x"142",x"040",x"9E6",x"9E5",x"9D5",x"AD5",x"AE4",x"AD5",x"140",x"040",x"7D5",x"6D4",x"6D4",x"7D4",x"AD4",x"AD4",x"AD4",x"AD5",x"140",x"140",x"140",x"140",x"00F",x"00F",x"00F",x"00B",x"234",x"240",x"AD5",x"AD5",x"BD6",x"BD6",x"AD5",x"AD5",x"140",x"140",x"8C5",x"8C5",x"8C5",x"8C5",x"AD6",x"AD5",x"BD6",x"BD6",x"140",x"141",x"143",x"134",x"00F",x"00F",x"00F",x"00B",x"647",x"652",x"AD6",x"BD6",x"651",x"551",x"8C5",x"7C4",x"AE6",x"AC6",x"551",x"652",x"652",x"552",x"240",x"240",x"552",x"552",x"240",x"132",x"018",x"00B",x"00F",x"00E",x"00C",x"109",x"646",x"652",x"AD7",x"AC6",x"552",x"552",x"9B6",x"9C6",x"BC6",x"CC7",x"742",x"743",x"742",x"652",x"240",x"240",x"553",x"553",x"230",x"234",x"00B",x"00F",x"00F",x"00C",x"53A",x"646",x"332",x"230",x"140",x"140",x"140",x"230",x"653",x"743",x"743",x"742",x"743",x"742",x"CC7",x"BC6",x"BD6",x"AD6",x"240",x"331",x"653",x"647",x"10B",x"00F",x"10C",x"209",x"636",x"743",x"330",x"340",x"230",x"240",x"240",x"330",x"743",x"833",x"833",x"833",x"844",x"742",x"CC7",x"CC6",x"CC6",x"BC7",x"230",x"330",x"643",x"636",x"208",x"10B",x"637",x"636",x"A66",x"A65",x"A64",x"964",x"752",x"642",x"964",x"964",x"A63",x"B64",x"A64",x"A64",x"833",x"733",x"743",x"743",x"642",x"642",x"643",x"743",x"A65",x"A66",x"736",x"737",x"843",x"843",x"A65",x"A64",x"B64",x"B65",x"832",x"843",x"B65",x"B64",x"A64",x"A63",x"A63",x"A64",x"832",x"943",x"833",x"833",x"843",x"843",x"833",x"843",x"A65",x"A65",x"833",x"833",x"A64",x"A64",x"743",x"843",x"833",x"843",x"733",x"843",x"833",x"843",x"732",x"742",x"B74",x"A63",x"B64",x"B54",x"B64",x"A64",x"A64",x"A65",x"833",x"834",x"843",x"833",x"A65",x"A64",x"A63",x"A64",x"843",x"743",x"834",x"834",x"844",x"844",x"834",x"834",x"844",x"743",x"A64",x"A63",x"B63",x"B64",x"A63",x"B63",x"B64",x"B64",x"833",x"834",x"834",x"843",x"A64",x"A63");
		-- Se define el mapa de bits para los arbustos del fondo
		constant arbusto : rom_cosas := ( x"00F",x"00F",x"00F",x"00C",x"004",x"000",x"000",x"000",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"000",x"000",x"000",x"003",x"00C",x"00F",x"00F",x"00F",x"00F",x"00F",x"00F",x"00E",x"00D",x"009",x"001",x"000",x"000",x"000",x"000",x"001",x"019",x"00C",x"00C",x"009",x"001",x"000",x"000",x"000",x"000",x"002",x"109",x"00C",x"00C",x"00D",x"00E",x"00F",x"00F",x"00D",x"006",x"001",x"BC8",x"BC6",x"BD6",x"BD6",x"BD6",x"BC9",x"001",x"003",x"003",x"001",x"8C8",x"8C5",x"AD6",x"AD7",x"140",x"142",x"002",x"003",x"003",x"006",x"00D",x"00F",x"00F",x"00C",x"003",x"000",x"BD7",x"AD5",x"BD6",x"BD6",x"AD6",x"AD7",x"010",x"000",x"000",x"010",x"8B6",x"8C6",x"BD7",x"AD7",x"150",x"040",x"000",x"000",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"230",x"240",x"000",x"000",x"140",x"140",x"140",x"140",x"8C6",x"8C6",x"010",x"000",x"000",x"000",x"8C5",x"8C4",x"AD6",x"BC8",x"000",x"003",x"00C",x"00F",x"00C",x"019",x"001",x"000",x"240",x"240",x"010",x"010",x"140",x"140",x"040",x"040",x"8C5",x"8B5",x"010",x"000",x"000",x"010",x"8C5",x"8C5",x"AD6",x"BD7",x"000",x"001",x"019",x"00C",x"003",x"001",x"AD8",x"AD6",x"BD5",x"BD5",x"AD5",x"AD6",x"140",x"040",x"7D6",x"7C6",x"010",x"010",x"AC6",x"AD6",x"BD6",x"AC7",x"010",x"010",x"140",x"140",x"AD6",x"BC8",x"001",x"003",x"000",x"000",x"AC7",x"AD6",x"BD6",x"BD5",x"AD5",x"AD5",x"150",x"050",x"7C5",x"7C6",x"010",x"010",x"AD6",x"AE5",x"AD5",x"BD7",x"000",x"010",x"140",x"140",x"AD6",x"BD7",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"AD6",x"AD5",x"AD5",x"AD6",x"040",x"050",x"7C5",x"7D5",x"7D4",x"7C5",x"010",x"000",x"8C6",x"7C5",x"AD6",x"AD7",x"000",x"000",x"000",x"000",x"003",x"002",x"001",x"000",x"000",x"010",x"AC7",x"AD6",x"9D5",x"AD6",x"140",x"040",x"7D4",x"6D4",x"6D4",x"7D5",x"010",x"000",x"8C6",x"7C5",x"AD6",x"BC8",x"000",x"001",x"002",x"003",x"00C",x"119",x"002",x"000",x"8C7",x"8C6",x"010",x"010",x"8C5",x"8C4",x"AD5",x"AD6",x"7D5",x"6D4",x"6D4",x"6D4",x"140",x"140",x"040",x"040",x"000",x"000",x"000",x"003",x"109",x"00C",x"00F",x"00B",x"003",x"000",x"7C5",x"7C5",x"010",x"010",x"7C5",x"8C5",x"AD5",x"AD6",x"7C5",x"6C5",x"6D4",x"7D4",x"050",x"050",x"050",x"150",x"010",x"000",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"7D6",x"6D4",x"7C4",x"7C5",x"040",x"140",x"140",x"040",x"150",x"050",x"050",x"050",x"6D5",x"6D5",x"6D5",x"6C5",x"140",x"241",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"7C5",x"6D3",x"6D3",x"7D4",x"050",x"140",x"040",x"141",x"040",x"140",x"141",x"040",x"6D5",x"6D4",x"6D4",x"6D4",x"040",x"140",x"000",x"001",x"019",x"00C",x"00F",x"00C",x"003",x"000",x"AD6",x"9E5",x"6D4",x"6D4",x"7D4",x"7C6",x"010",x"000",x"000",x"000",x"000",x"010",x"7C5",x"6D4",x"6D3",x"7D4",x"AE6",x"BD6",x"BD6",x"BC8",x"001",x"003",x"00C",x"009",x"001",x"010",x"AD6",x"9E5",x"6D4",x"6D4",x"7C5",x"7C6",x"010",x"000",x"000",x"000",x"000",x"000",x"8C6",x"7C5",x"7D4",x"7D4",x"9D5",x"AD5",x"AD4",x"BD6",x"000",x"000",x"003",x"001",x"8C7",x"7D5",x"7C4",x"7D4",x"6D4",x"6D5",x"010",x"010",x"8C6",x"7C5",x"7C5",x"8C5",x"AD6",x"BC7",x"000",x"010",x"7C5",x"7D4",x"040",x"140",x"7C4",x"8C5",x"000",x"001",x"003",x"001",x"7B6",x"7C5",x"8C5",x"7C5",x"6D4",x"6C4",x"010",x"010",x"8C6",x"8D6",x"6C5",x"7D4",x"AD5",x"AD6",x"000",x"010",x"7C5",x"7D5",x"150",x"040",x"7C6",x"7C7",x"002",x"004",x"00C",x"009",x"001",x"000",x"000",x"010",x"9D5",x"9E5",x"7C5",x"8C6",x"000",x"000",x"140",x"040",x"140",x"140",x"AD6",x"9D5",x"6D4",x"6C5",x"040",x"140",x"010",x"001",x"019",x"00C",x"00F",x"00C",x"003",x"000",x"000",x"000",x"AD6",x"9D5",x"7C4",x"7D6",x"010",x"010",x"140",x"040",x"040",x"040",x"AD6",x"9D5",x"7D5",x"7D6",x"140",x"240",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"241",x"140",x"140",x"040",x"6D5",x"6D4",x"7D5",x"7C6",x"040",x"140",x"140",x"140",x"140",x"140",x"040",x"050",x"AD6",x"AC6",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"130",x"140",x"241",x"140",x"7C6",x"7C5",x"7C5",x"7C6",x"140",x"140",x"141",x"141",x"241",x"130",x"141",x"140",x"AD7",x"BC7",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"010",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"003",x"00C",x"00F",x"00F",x"00C",x"003",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"003",x"10C",x"00F");
		
		-- Matriz para manejar un diseño del fondo
		type rom_cosas2 is array (0 to 1599) of std_logic_vector(11 downto 0);
		-- Se define el mapa de bits para las lunas del fondo
		constant luna : rom_cosas2 := ( x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2E2",x"595",x"787",x"788",x"788",x"778",x"778",x"887",x"887",x"878",x"888",x"787",x"787",x"888",x"878",x"878",x"595",x"1E2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E2",x"2E2",x"2E2",x"4D4",x"695",x"887",x"787",x"778",x"888",x"888",x"777",x"887",x"778",x"788",x"887",x"787",x"877",x"878",x"878",x"696",x"3D4",x"1E2",x"1E2",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2E2",x"4A4",x"696",x"595",x"696",x"565",x"655",x"555",x"666",x"555",x"555",x"666",x"555",x"BCC",x"BCC",x"BBB",x"BCB",x"CCC",x"CBC",x"878",x"777",x"696",x"595",x"595",x"4A4",x"2E2",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"2E1",x"2E2",x"2E2",x"4D4",x"696",x"888",x"878",x"777",x"655",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"BCC",x"BCC",x"BCB",x"CCB",x"BBC",x"CCC",x"888",x"877",x"887",x"787",x"777",x"696",x"4D4",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"4A3",x"595",x"595",x"696",x"565",x"555",x"555",x"565",x"555",x"565",x"656",x"655",x"655",x"665",x"655",x"656",x"555",x"555",x"CCC",x"BBC",x"BBC",x"BCC",x"BCB",x"BCB",x"CBB",x"CBC",x"878",x"787",x"696",x"3B3",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"3D4",x"696",x"877",x"777",x"788",x"565",x"555",x"555",x"555",x"565",x"555",x"655",x"655",x"554",x"665",x"555",x"555",x"656",x"656",x"BBC",x"CCC",x"CCC",x"BBB",x"BCB",x"CCB",x"CBC",x"CBC",x"878",x"777",x"778",x"696",x"4D3",x"1E1",x"1F0",x"0F0",x"0F0",x"0F0",x"0F1",x"1E2",x"3A4",x"696",x"787",x"878",x"666",x"555",x"555",x"555",x"565",x"565",x"555",x"555",x"555",x"555",x"CCB",x"BBB",x"BCB",x"BCB",x"555",x"556",x"566",x"556",x"CBB",x"CCB",x"CBB",x"CCB",x"CBB",x"CBC",x"BCB",x"CCC",x"888",x"787",x"696",x"4A4",x"2E1",x"0F0",x"0F0",x"0F0",x"0F0",x"2E3",x"596",x"878",x"888",x"878",x"556",x"555",x"555",x"555",x"555",x"565",x"555",x"566",x"555",x"555",x"CCC",x"CBC",x"BCB",x"BCB",x"555",x"666",x"555",x"566",x"CCB",x"CBB",x"CBC",x"CCC",x"BBC",x"BBC",x"BCC",x"BBB",x"888",x"778",x"888",x"595",x"2E2",x"0F0",x"0F0",x"0F0",x"0F0",x"2E2",x"595",x"877",x"655",x"555",x"556",x"556",x"BBC",x"CCC",x"555",x"565",x"556",x"556",x"555",x"555",x"556",x"556",x"555",x"665",x"555",x"556",x"566",x"555",x"655",x"555",x"CCC",x"CCC",x"BBC",x"CCC",x"BBC",x"CCC",x"CCC",x"BBB",x"787",x"595",x"2E1",x"0F0",x"0F0",x"0F0",x"2E2",x"4D4",x"696",x"877",x"655",x"555",x"556",x"556",x"CCC",x"BBB",x"666",x"555",x"556",x"556",x"556",x"556",x"666",x"556",x"555",x"555",x"555",x"556",x"555",x"555",x"555",x"666",x"BBB",x"CCC",x"BBC",x"BBC",x"CCC",x"CCC",x"CCC",x"CCC",x"787",x"595",x"3D3",x"1E1",x"0F0",x"0F0",x"595",x"595",x"564",x"655",x"555",x"555",x"655",x"655",x"656",x"666",x"556",x"556",x"656",x"655",x"555",x"566",x"555",x"555",x"665",x"665",x"555",x"555",x"556",x"555",x"555",x"555",x"565",x"555",x"CCC",x"CCC",x"CCB",x"BBB",x"BBB",x"BBB",x"778",x"787",x"696",x"3A4",x"2E2",x"0F0",x"888",x"887",x"555",x"555",x"555",x"555",x"655",x"655",x"656",x"555",x"666",x"555",x"655",x"655",x"555",x"556",x"555",x"665",x"555",x"555",x"555",x"555",x"556",x"555",x"555",x"665",x"565",x"555",x"CCC",x"BBB",x"BBB",x"BCB",x"CCC",x"BBC",x"888",x"878",x"878",x"696",x"4C4",x"3E3",x"776",x"887",x"555",x"555",x"566",x"556",x"555",x"555",x"666",x"555",x"555",x"655",x"655",x"656",x"556",x"555",x"655",x"655",x"555",x"555",x"655",x"555",x"666",x"555",x"555",x"565",x"555",x"656",x"000",x"000",x"CCC",x"CCC",x"CBC",x"CBC",x"CBC",x"CBC",x"878",x"777",x"696",x"595",x"887",x"877",x"555",x"556",x"555",x"555",x"665",x"555",x"556",x"555",x"655",x"665",x"555",x"555",x"566",x"556",x"655",x"656",x"555",x"555",x"655",x"655",x"555",x"566",x"555",x"555",x"555",x"556",x"000",x"000",x"CBC",x"BBC",x"CBC",x"CBB",x"CBB",x"CBB",x"878",x"878",x"788",x"787",x"777",x"888",x"555",x"656",x"CCC",x"BCB",x"555",x"556",x"555",x"555",x"555",x"655",x"655",x"555",x"555",x"555",x"556",x"555",x"BBB",x"CCC",x"555",x"555",x"666",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"BBB",x"CCC",x"CCC",x"BBC",x"CCB",x"CCB",x"777",x"777",x"887",x"787",x"888",x"778",x"556",x"665",x"BBB",x"CCB",x"655",x"656",x"556",x"556",x"655",x"555",x"655",x"555",x"565",x"566",x"566",x"566",x"BCC",x"BCC",x"555",x"666",x"555",x"565",x"000",x"000",x"000",x"000",x"000",x"000",x"CCB",x"BCB",x"BBB",x"CCC",x"BBB",x"BBB",x"887",x"787",x"787",x"787",x"888",x"778",x"556",x"555",x"554",x"655",x"655",x"556",x"556",x"556",x"BCC",x"CCB",x"000",x"000",x"566",x"555",x"555",x"555",x"565",x"555",x"CCC",x"CCC",x"CCC",x"BCC",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"BBB",x"BBB",x"BBB",x"CCB",x"CBB",x"CBB",x"CCB",x"CCB",x"777",x"788",x"778",x"778",x"555",x"565",x"655",x"554",x"665",x"556",x"556",x"556",x"BCC",x"CCB",x"000",x"000",x"555",x"566",x"556",x"666",x"555",x"555",x"BBB",x"BBB",x"BBB",x"CCC",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"CCC",x"CCC",x"CCB",x"BBB",x"CBC",x"CCC",x"BBB",x"CCB",x"888",x"778",x"887",x"887",x"CBB",x"CBB",x"655",x"555",x"000",x"000",x"665",x"555",x"BCB",x"CCB",x"655",x"555",x"566",x"555",x"555",x"555",x"BBB",x"CCC",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"BBB",x"BBB",x"CCC",x"BBB",x"000",x"000",x"CCC",x"CBC",x"CCC",x"CCB",x"887",x"777",x"887",x"777",x"CCC",x"CBB",x"656",x"555",x"000",x"000",x"555",x"655",x"CCB",x"BBB",x"665",x"555",x"555",x"555",x"555",x"666",x"BBB",x"CCC",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"BBB",x"CCC",x"000",x"000",x"BBC",x"CBC",x"BBB",x"BBB",x"888",x"887",x"778",x"778",x"788",x"788",x"555",x"655",x"000",x"000",x"655",x"555",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"CCC",x"BBB",x"BBB",x"CCC",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"BBB",x"BBB",x"CCC",x"BBB",x"CCB",x"CCB",x"000",x"000",x"BCB",x"CCC",x"777",x"777",x"888",x"788",x"788",x"788",x"555",x"656",x"000",x"000",x"666",x"555",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"CCC",x"CCC",x"BBB",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"BBB",x"CCB",x"CBB",x"CCB",x"000",x"000",x"CCB",x"BCC",x"888",x"788",x"787",x"787",x"787",x"777",x"656",x"556",x"556",x"566",x"555",x"555",x"FFF",x"FFF",x"FFF",x"FFF",x"BBB",x"BCC",x"CCC",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"FFF",x"FFF",x"BBB",x"CCC",x"BBB",x"BBB",x"CCC",x"CCC",x"BBB",x"CCC",x"CCC",x"BCC",x"BBC",x"BBC",x"778",x"888",x"787",x"887",x"777",x"787",x"666",x"556",x"566",x"556",x"565",x"565",x"FFF",x"FFF",x"FFF",x"FFF",x"BCC",x"BCC",x"CCC",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"FFF",x"FFF",x"CCC",x"CCC",x"CCC",x"CCC",x"CCC",x"BCB",x"BCB",x"BCC",x"BBC",x"CCC",x"BCC",x"CCC",x"888",x"778",x"878",x"878",x"888",x"888",x"000",x"000",x"555",x"655",x"CCB",x"CCB",x"FFF",x"FFF",x"BCC",x"BCB",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"BBB",x"BBB",x"CCC",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"BBB",x"CCC",x"BBB",x"CCC",x"BCB",x"BCC",x"CBC",x"CBC",x"CCC",x"BCB",x"788",x"788",x"878",x"878",x"878",x"777",x"000",x"000",x"655",x"655",x"CBB",x"CBB",x"FFF",x"FFF",x"BBB",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"BBB",x"CCC",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"BBB",x"CCC",x"BBB",x"CCB",x"BBB",x"CBC",x"CBC",x"BCC",x"BCC",x"778",x"778",x"878",x"988",x"878",x"888",x"BCB",x"BCB",x"655",x"655",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"BBB",x"CCC",x"000",x"000",x"FFF",x"FFF",x"CCC",x"CCC",x"BBB",x"CCC",x"CCC",x"CCC",x"BBB",x"CCC",x"CBB",x"CBB",x"CCC",x"BBB",x"878",x"878",x"595",x"685",x"787",x"888",x"BBB",x"BCB",x"655",x"555",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"CCC",x"BBB",x"000",x"000",x"FFF",x"FFF",x"BBB",x"BBB",x"CCC",x"CCC",x"CCC",x"BBB",x"BCB",x"BBB",x"CCB",x"CBB",x"BBB",x"BBC",x"878",x"878",x"1E2",x"3D4",x"696",x"777",x"CCB",x"CCC",x"555",x"556",x"566",x"556",x"666",x"555",x"556",x"555",x"555",x"555",x"FFF",x"FFF",x"BBB",x"BBB",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"CCC",x"BBB",x"CCC",x"CCC",x"BCB",x"BCB",x"BCB",x"CCC",x"888",x"878",x"888",x"777",x"0F0",x"1E2",x"5A5",x"887",x"CBB",x"CBC",x"656",x"556",x"556",x"556",x"555",x"555",x"656",x"556",x"665",x"555",x"FFF",x"FFF",x"CCC",x"CCC",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"BBB",x"CCC",x"CCC",x"BBB",x"CCC",x"BCB",x"BCB",x"BCC",x"BCC",x"878",x"787",x"696",x"5A5",x"0F0",x"2E2",x"595",x"888",x"878",x"888",x"BCB",x"BCB",x"555",x"556",x"555",x"665",x"556",x"556",x"555",x"665",x"FFF",x"FFF",x"BBB",x"CCC",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"BBB",x"CCC",x"BBB",x"CCC",x"CCC",x"BBB",x"CBB",x"CBB",x"788",x"888",x"877",x"696",x"4D4",x"2E2",x"0F0",x"1E2",x"4A3",x"696",x"787",x"778",x"CCB",x"CCC",x"556",x"556",x"555",x"555",x"655",x"655",x"555",x"555",x"FFF",x"FFF",x"CCC",x"BBB",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"CCC",x"CCC",x"BBB",x"CCC",x"CCC",x"BBB",x"CCC",x"CBB",x"CBB",x"888",x"777",x"887",x"595",x"2E2",x"0F0",x"0F0",x"0F0",x"1E1",x"4C4",x"696",x"787",x"CCB",x"CBB",x"556",x"556",x"565",x"555",x"555",x"655",x"555",x"565",x"FFF",x"FFF",x"000",x"000",x"FFF",x"FFF",x"000",x"000",x"CCC",x"BBB",x"CCC",x"BBB",x"CCC",x"BBB",x"000",x"000",x"777",x"887",x"777",x"888",x"888",x"595",x"2E3",x"0F1",x"0F0",x"0F0",x"0F0",x"2E2",x"595",x"887",x"CBB",x"CBC",x"556",x"556",x"565",x"666",x"555",x"665",x"555",x"555",x"FFF",x"FFF",x"000",x"000",x"FFF",x"FFF",x"000",x"000",x"BBB",x"BBB",x"CCC",x"CCC",x"CCC",x"CCC",x"000",x"000",x"887",x"888",x"877",x"787",x"696",x"3A4",x"2E2",x"0F1",x"0F0",x"0F0",x"0F0",x"2E2",x"5A5",x"777",x"988",x"878",x"CBC",x"CCC",x"BBB",x"BCB",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"BBB",x"CCC",x"BBB",x"CCC",x"BBB",x"000",x"000",x"888",x"888",x"777",x"878",x"878",x"696",x"4D4",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"3A3",x"696",x"787",x"878",x"CBC",x"CBC",x"CCC",x"CCC",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"CCC",x"BBB",x"CCC",x"CCC",x"CCC",x"BBB",x"000",x"000",x"777",x"888",x"887",x"787",x"696",x"4A4",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"4C3",x"696",x"888",x"878",x"878",x"BBB",x"BCB",x"BBB",x"CCC",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"BBB",x"CCC",x"BBB",x"BBB",x"000",x"000",x"777",x"777",x"888",x"888",x"888",x"696",x"4D4",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"3B3",x"596",x"787",x"888",x"CCC",x"BCB",x"CCB",x"CCB",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"CCC",x"BBB",x"CCC",x"CCC",x"000",x"000",x"777",x"888",x"777",x"787",x"696",x"3A4",x"1E1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"3D3",x"696",x"778",x"788",x"777",x"777",x"887",x"BBB",x"CCB",x"FFF",x"FFF",x"FFF",x"FFF",x"888",x"777",x"777",x"888",x"777",x"888",x"888",x"777",x"888",x"777",x"777",x"696",x"4C5",x"2E2",x"0F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"1E1",x"595",x"788",x"778",x"888",x"878",x"887",x"CCB",x"BCB",x"FFF",x"FFF",x"FFF",x"FFF",x"777",x"777",x"888",x"777",x"888",x"777",x"888",x"888",x"777",x"888",x"888",x"596",x"2D3",x"0F1",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");
		
		-- Matriz para manejar las vidas del juego
		type rom_vida is array (0 to 623) of std_logic_vector(11 downto 0);
		-- Se define el mapa de bits para el corazón
		constant vida : rom_vida := ( x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"000",x"000",x"000",x"000",x"000",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"000",x"000",x"000",x"000",x"000",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"FFE",x"200",x"200",x"200",x"200",x"200",x"100",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"200",x"200",x"200",x"200",x"200",x"200",x"0F0",x"0F0",x"0F0",x"0F0",x"FEF",x"0F0",x"000",x"200",x"A21",x"C11",x"C10",x"D11",x"D11",x"B22",x"200",x"000",x"0F0",x"0F0",x"000",x"200",x"B22",x"C11",x"D11",x"C10",x"D11",x"B21",x"200",x"000",x"0F0",x"0F0",x"0F0",x"FEF",x"100",x"400",x"B11",x"C10",x"D11",x"D00",x"F00",x"D00",x"500",x"200",x"0F0",x"FEE",x"200",x"400",x"D11",x"F00",x"F00",x"F00",x"F00",x"D00",x"500",x"200",x"0F0",x"0F0",x"000",x"200",x"A21",x"B11",x"FED",x"FEE",x"FEE",x"FED",x"D11",x"F00",x"D11",x"A21",x"200",x"200",x"A11",x"D10",x"E00",x"F00",x"F00",x"F00",x"F00",x"E00",x"D00",x"B22",x"200",x"000",x"000",x"200",x"D11",x"C10",x"FEE",x"0F0",x"FFE",x"FED",x"D01",x"F00",x"F00",x"D10",x"400",x"400",x"D11",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"C11",x"200",x"000",x"000",x"200",x"C11",x"C11",x"FEF",x"FEF",x"B22",x"D11",x"E00",x"F00",x"F00",x"E00",x"D10",x"D11",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D11",x"200",x"000",x"000",x"200",x"D11",x"D01",x"FDE",x"FDE",x"D00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D11",x"200",x"000",x"000",x"300",x"D10",x"F00",x"D01",x"D01",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D11",x"300",x"000",x"000",x"300",x"D11",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D10",x"300",x"000",x"000",x"200",x"C10",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"C10",x"200",x"000",x"000",x"100",x"A21",x"D10",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"E00",x"D00",x"A22",x"100",x"000",x"0F0",x"0F0",x"200",x"400",x"D11",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D01",x"400",x"100",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"100",x"A12",x"D01",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D01",x"B22",x"200",x"000",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"200",x"500",x"D00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D00",x"400",x"200",x"FEE",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"200",x"B22",x"D01",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"E00",x"D01",x"B22",x"200",x"000",x"0F0",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"FEE",x"200",x"400",x"E11",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D01",x"400",x"200",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"100",x"A11",x"D10",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"D01",x"A22",x"200",x"000",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"EFF",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"0F0",x"0F0",x"200",x"400",x"D00",x"F00",x"F00",x"F00",x"F00",x"D11",x"400",x"200",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"EFF",x"EFF",x"0F0",x"0F0",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"200",x"A22",x"D10",x"F00",x"E00",x"D11",x"A22",x"100",x"000",x"FFE",x"FFE",x"0F0",x"FEF",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"100",x"400",x"E11",x"D00",x"500",x"200",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"000",x"200",x"B21",x"B21",x"200",x"000",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"EFF",x"0F0",x"0F0",x"0F0",x"FFE",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"FFE",x"200",x"200",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"EFF",x"0F0",x"EFF",x"0F0",x"FFE",x"FFE",x"FFE",x"0F0",x"0F0",x"0F0",x"FFE",x"FFE",x"000",x"000",x"EFF",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0",x"0F0");

	begin 
		-- Las siguiente lineas se encargan de dibujar la sección de datos
		if(xcur>160+540 and xcur<=160+640 and ycur>45 and ycur<=45+480) then
			-- Margen izquierdo
			if(xcur>160+540 and xcur<=160+550) then
				pos_dx := ((160+550) - xcur);
				for y in 0 to 48 loop
					pos_dy := ((45+(y*10)+10) - ycur);
					exit when (ycur>(45+(y*10)) and ycur<=(45+(y*10)+10)); 
				end loop;
				
				if(margen_v(pos_dy)(pos_dx) = '1') then
					rgb <= x"f04";
				else
					rgb <= x"000";
				end if;
			-- Margen derecho
			elsif(xcur>160+630 and xcur<=160+640) then
				pos_dx := ((160+640) - xcur);
				for y in 0 to 48 loop
					pos_dy := ((45+(y*10)+10) - ycur);
					exit when (ycur>(45+(y*10)) and ycur<=(45+(y*10)+10)); 
				end loop;
				
				if(margen_v(pos_dy)(pos_dx) = '1') then
					rgb <= x"f04";
				else
					rgb <= x"000";
				end if;
			-- Margen superior
			elsif(xcur>160+550 and xcur<=160+630) then
				if (ycur>45 and ycur<=45+10) then
					pos_dy := ((45+10)-ycur);
					
					for x in 55 to 64 loop
						pos_dx := ((160+(x*10)+10) - xcur);
						exit when (xcur>(160+(x*10)) and xcur<=(160+(x*10)+10)); 
					end loop;
					
					if(margen_h(pos_dy)(pos_dx) = '1') then
						rgb <= x"f04";
					else
						rgb <= x"000";
					end if;
				-- La siguiente sección se dedica a dibujar los corazones de la vida
				elsif(ycur>45+15 and ycur<=45+39) then
					if(life > 0) then
						pos_dy := (24-((45+39)-ycur));
						
						if(life = 3) then
							if(xcur>160+551 and xcur<=160+577) then
								pos_dx := (26-((160+577)-xcur));
								al := 1;
							elsif(xcur>160+577 and xcur<=160+603) then
								pos_dx := (26-((160+603)-xcur));
								al := 1;
							elsif(xcur>160+603 and xcur<=160+629) then
								pos_dx := (26-((160+629)-xcur));
								al := 1;
							else
								al := 0;
							end if;
						elsif(life = 2) then
							if(xcur>160+551 and xcur<=160+577) then
								pos_dx := (26-((160+577)-xcur));
								al := 1;
							elsif(xcur>160+577 and xcur<=160+603) then
								pos_dx := (26-((160+603)-xcur));
								al := 1;
							else
								al := 0;
							end if;
						elsif(life = 1) then
							if(xcur>160+551 and xcur<=160+577) then
								pos_dx := (26-((160+577)-xcur));
								al := 1;
							else
								al := 0;
							end if;
						end if;
						
						if (al = 1) then
							if (vida(pos_dx + (26*pos_dy)) /= x"0f0") then
								rgb <= vida(pos_dx + (26*pos_dy));
							else 
								rgb <= x"000";
							end if;
						else
							rgb <= x"000";
						end if;
					else
						rgb <= x"000";
					end if;
				-- Letrero score
				elsif (ycur>45+100 and ycur<=45+115) then
					if (xcur>160+553 and xcur<=160+628) then
						pos_dx := (74-((160+628) - xcur));
						pos_dy := (14-((45+115)-ycur));
						
						if(l_score(pos_dy)(pos_dx) = '1') then
							rgb <= x"fff";
						else
							rgb <= x"000";
						end if;
					else
						rgb <= x"000";
					end if;
				-- Letrero nivel
				elsif (ycur>45+200 and ycur<=45+215) then
					if (xcur>160+553 and xcur<=160+628) then
						pos_dx := (74-((160+628) - xcur));
						pos_dy := (14-((45+215)-ycur));
						
						if(l_nivel(pos_dy)(pos_dx) = '1') then
							rgb <= x"fff";
						else
							rgb <= x"000";
						end if;
					else
						rgb <= x"000";
					end if;
				elsif (ycur>45+120 and ycur<=45+135) then
					pos_dy := (14-((45+135)-ycur));
					-- Score millares
					if (xcur>160+550 and xcur<=160+565) then
						pos_dx := (14-((160+565) - xcur));
						if(sc_mm = 0) then
							if(cero(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 1) then
							if(uno(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 2) then
							if(dos(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 3) then
							if(tres(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 4) then
							if(cuatro(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 5) then
							if(cinco(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 6) then
							if(seis(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 7) then
							if(siete(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 8) then
							if(ocho(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_mm = 9) then
							if(nueve(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					-- Score miles
					elsif (xcur>160+566 and xcur<=160+581) then
						pos_dx := (14-((160+581) - xcur));
						if(sc_m = 0) then
							if(cero(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 1) then
							if(uno(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 2) then
							if(dos(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 3) then
							if(tres(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 4) then
							if(cuatro(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 5) then
							if(cinco(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 6) then
							if(seis(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 7) then
							if(siete(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 8) then
							if(ocho(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_m = 9) then
							if(nueve(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					-- Score centenas
					elsif (xcur>160+582 and xcur<=160+597) then
						pos_dx := (14-((160+597) - xcur));
						if(sc_c = 0) then
							if(cero(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 1) then
							if(uno(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 2) then
							if(dos(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 3) then
							if(tres(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 4) then
							if(cuatro(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 5) then
							if(cinco(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 6) then
							if(seis(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 7) then
							if(siete(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 8) then
							if(ocho(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_c = 9) then
							if(nueve(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					-- Score decenas
					elsif (xcur>160+598 and xcur<=160+613) then
						pos_dx := (14-((160+613) - xcur));
						if(sc_d = 0) then
							if(cero(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 1) then
							if(uno(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 2) then
							if(dos(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 3) then
							if(tres(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 4) then
							if(cuatro(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 5) then
							if(cinco(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 6) then
							if(seis(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 7) then
							if(siete(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 8) then
							if(ocho(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(sc_d = 9) then
							if(nueve(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					-- Score unidades
					elsif (xcur>160+614 and xcur<=160+629) then
						pos_dx := (14-((160+629) - xcur));
						if(sc_u = 0) then
							if(cero(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					else
						rgb <= x"000";
					end if;
				-- Número nivel
				elsif (ycur>45+220 and ycur<=45+235) then
					if (xcur>160+582 and xcur<=160+597) then
						pos_dx := (14-((160+597) - xcur));
						pos_dy := (14-((45+235)-ycur));
						
						if(nivel = 1) then
							if(uno(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(nivel = 2) then
							if(dos(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(nivel = 3) then
							if(tres(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						elsif(nivel = 4) then
							if(cuatro(pos_dy)(pos_dx) = '1') then
								rgb <= x"fff";
							else
								rgb <= x"000";
							end if;
						end if;
					else
						rgb <= x"000";
					end if;
				-- Margen inferior
				elsif (ycur>45+470 and ycur<=45+480) then
					pos_dy := ((45+480)-ycur);
					
					for x in 55 to 64 loop
						pos_dx := ((160+(x*10)+10) - xcur);
						exit when (xcur>(160+(x*10)) and xcur<=(160+(x*10)+10)); 
					end loop;
					
					if(margen_h(pos_dy)(pos_dx) = '1') then
						rgb <= x"f04";
					else
						rgb <= x"000";
					end if;
				else
					rgb <= x"000";
				end if;
			end if;
		-- Las siguientes líneas se dedican a dibujar la sección del juego
		elsif (nivel = 1 or nivel = 2) then
			-- Fondo verde izquierdo, nivel 1 arbustos y nivel 2 flores
			if(xcur>160+120 and xcur<=160+210 and ycur>45 and ycur<=45+480) then
				if (xcur>160+120+10 and xcur<=160+120+36 and ycur>45+10 and ycur<=45+34) then
					pos_dx := (25-((160+120+36) - xcur));
					pos_dy := (23-((45+34) - ycur));
					ac := 1;
				elsif (xcur>160+120+54 and xcur<=160+120+80 and ycur>45+100 and ycur<=45+124) then
					pos_dx := (25-((160+120+80) - xcur));
					pos_dy := (23-((45+124) - ycur));
					ac := 1;
				elsif (xcur>160+120+10 and xcur<=160+120+36 and ycur>45+200 and ycur<=45+224) then
					pos_dx := (25-((160+120+36) - xcur));
					pos_dy := (23-((45+224) - ycur));
					ac := 1;
				elsif (xcur>160+120+54 and xcur<=160+120+80 and ycur>45+300 and ycur<=45+324) then
					pos_dx := (25-((160+120+80) - xcur));
					pos_dy := (23-((45+324) - ycur));
					ac := 1;	
				elsif (xcur>160+120+10 and xcur<=160+120+36 and ycur>45+400 and ycur<=45+424) then
					pos_dx := (25-((160+120+36) - xcur));
					pos_dy := (23-((45+424) - ycur));
					ac := 1;
				else
					ac := 0;
				end if;
				
				if (ac = 0) then
					if(nivel = 1) then
						rgb <= x"bf0";
					elsif (nivel = 2) then
						rgb <= x"8f0";
					end if;
				elsif(nivel = 1) then					
					if (arbusto(pos_dx + (26*pos_dy)) /= x"00f") then
						rgb <= arbusto(pos_dx + (26*pos_dy));
					else 
						rgb <= x"bf0";
					end if;
				elsif (nivel = 2) then
					if (flores(pos_dx + (26*pos_dy)) /= x"00f") then
						rgb <= flores(pos_dx + (26*pos_dy));
					else 
						rgb <= x"8f0";
					end if;
				end if;
			-- Fondo verde derecho, nivel 1 arbustos y nivel 2 flores
			elsif(xcur>160+330 and xcur<=160+420 and ycur>45 and ycur<=45+480) then
				if (xcur>160+330+10 and xcur<=160+330+36 and ycur>45+10 and ycur<=45+34) then
					pos_dx := (25-((160+330+36) - xcur));
					pos_dy := (23-((45+34) - ycur));
					ac := 1;
				elsif (xcur>160+330+54 and xcur<=160+330+80 and ycur>45+100 and ycur<=45+124) then
					pos_dx := (25-((160+330+80) - xcur));
					pos_dy := (23-((45+124) - ycur));
					ac := 1;
				elsif (xcur>160+330+10 and xcur<=160+330+36 and ycur>45+200 and ycur<=45+224) then
					pos_dx := (25-((160+330+36) - xcur));
					pos_dy := (23-((45+224) - ycur));
					ac := 1;
				elsif (xcur>160+330+54 and xcur<=160+330+80 and ycur>45+300 and ycur<=45+324) then
					pos_dx := (25-((160+330+80) - xcur));
					pos_dy := (23-((45+324) - ycur));	
					ac := 1;	
				elsif (xcur>160+330+10 and xcur<=160+330+36 and ycur>45+400 and ycur<=45+424) then
					pos_dx := (25-((160+330+36) - xcur));
					pos_dy := (23-((45+424) - ycur));
					ac := 1;
				else
					ac := 0;
				end if;
				
				if (ac = 0) then
					if(nivel = 1) then
						rgb <= x"bf0";
					elsif (nivel = 2) then
						rgb <= x"8f0";
					end if;
				elsif(nivel = 1) then					
					if (arbusto(pos_dx + (26*pos_dy)) /= x"00f") then
						rgb <= arbusto(pos_dx + (26*pos_dy));
					else 
						rgb <= x"bf0";
					end if;
				elsif (nivel = 2) then
					if (flores(pos_dx + (26*pos_dy)) /= x"00f") then
						rgb <= flores(pos_dx + (26*pos_dy));
					else 
						rgb <= x"8f0";
					end if;
				end if;
			-- Piso lado izquierdo
			elsif(xcur>160 and xcur<=160+120 and ycur>45 and ycur<=45+480) then
				pos_dx := (239-((160+120)-xcur));
					
				for y in 0 to 30 loop
					pos_dy := (15-((45+(y*16)+16) - ycur));
					exit when (ycur>(45+(y*16)) and ycur<=(45+(y*16)+16)); 
				end loop;
				
				if(nivel = 1) then
					rgb<= piso1(pos_dx + (120*pos_dy));
				elsif(nivel = 2) then
					rgb<= piso2(pos_dx + (120*pos_dy));
				end if;
			-- Piso centro
			elsif(xcur>160+210 and xcur<=160+330 and ycur>45 and ycur<=45+480) then
				pos_dx := (239-((160+330)-xcur));
					
				for y in 0 to 30 loop
					pos_dy := (15-((45+(y*16)+16) - ycur));
					exit when (ycur>(45+(y*16)) and ycur<=(45+(y*16)+16)); 
				end loop;
				
				if(nivel = 1) then
					rgb<= piso2(pos_dx + (120*pos_dy));
				elsif(nivel = 2) then
					rgb<= piso1(pos_dx + (120*pos_dy));
				end if;
			-- Piso lado derecho
			elsif(xcur>160+420 and xcur<=160+540 and ycur>45 and ycur<=45+480) then
				pos_dx := (239-((160+540)-xcur));
					
				for y in 0 to 30 loop
					pos_dy := (15-((45+(y*16)+16) - ycur));
					exit when (ycur>(45+(y*16)) and ycur<=(45+(y*16)+16)); 
				end loop;
				
				if(nivel = 1) then
					rgb<= piso1(pos_dx + (120*pos_dy));
				elsif(nivel = 2) then
					rgb<= piso2(pos_dx + (120*pos_dy));
				end if;
			end if;
		elsif (nivel = 3 or nivel = 4) then
			-- Fondo espacio 
			-- El nivel 3 solo es fondo negro con estrellas y en el nivel 4 hay lunas
			if(xcur>160 and xcur<=160+540 and ycur>45 and ycur<=45+480) then
				if (nivel = 4) then
					if (xcur>160+10 and xcur<=160+50 and ycur>45+10 and ycur<=45+50) then
						pos_dx := ((160+50) - xcur);
						pos_dy := ((45+50) - ycur);
						ae := 1;
					elsif (xcur>160+120+20 and xcur<=160+120+60 and ycur>45+300 and ycur<=45+340) then
						pos_dx := ((160+120+60) - xcur);
						pos_dy := ((45+340) - ycur);
						ae := 1;
					elsif (xcur>160+360+20 and xcur<=160+360+60 and ycur>45+80 and ycur<=45+120) then
						pos_dx := ((160+360+60) - xcur);
						pos_dy := ((45+120) - ycur);
						ae := 1;
					elsif (xcur>160+480+10 and xcur<=160+480+50 and ycur>45+420 and ycur<=45+460) then
						pos_dx := ((160+480+50) - xcur);
						pos_dy := ((45+460) - ycur);
						ae := 1;
					else
						ae := 0;
					end if;
					
					if (ae = 1) then
						if (luna(pos_dx + (40*pos_dy)) /= x"0f0") then
							rgb <= luna(pos_dx + (40*pos_dy));
						else 
							rgb <= x"222";
						end if;
					end if;
				else
					ae := 0;
				end if;
				
				if (ae = 0) then
					for y in 0 to 30 loop
						pos_dy := ((45+(y*16)+16) - ycur);
						ay := y;
						exit when (ycur>(45+(y*16)) and ycur<=(45+(y*16)+16)); 
					end loop;
						
					for x in 0 to 5 loop
						pos_dx := ((160+(x*120)+120) - xcur);
						ax := x;
						exit when (xcur>(160+(x*120)) and xcur<=(160+(x*120)+120)); 
					end loop;

					if (ay=0 or ay=3 or ay=6 or ay=9 or ay=12 or ay=15 or ay=18 or ay=21 or ay=24 or ay=27 or ay=30) then	
						if (ax = 0 or ax = 3) then
							rgb <= piso3(pos_dx + (120*pos_dy));
						elsif (ax = 1 or ax = 4) then
							rgb <= x"222";
						elsif (ax = 2 or ax = 5) then
							rgb <= piso4(pos_dx + (120*pos_dy));
						end if;
					elsif (ay=1 or ay=4 or ay=7 or ay=10 or ay=13 or ay=16 or ay=19 or ay=22 or ay=25 or ay=28) then
						if (ax = 0 or ax = 3) then
							rgb <= piso4(pos_dx + (120*pos_dy));
						elsif (ax = 1 or ax = 4) then
							rgb <= piso3(pos_dx + (120*pos_dy));
						elsif (ax = 2 or ax = 5) then
							rgb <= x"222";
						end if;
					elsif (ay=2 or ay=5 or ay=8 or ay=11 or ay=14 or ay=17 or ay=20 or ay=23 or ay=26 or ay=29) then
						if (ax = 0 or ax = 3) then
							rgb <= x"222";
						elsif (ax = 1 or ax = 4) then
							rgb <= piso4(pos_dx + (120*pos_dy));
						elsif (ax = 2 or ax = 5) then
							rgb <= piso3(pos_dx + (120*pos_dy));
						end if;	
					end if;
				end if;
			end if;
		end if;
	end background_play;
end background;